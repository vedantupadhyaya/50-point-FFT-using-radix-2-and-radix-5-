/////////////////////RADIX-2 ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module radix_2(clk,re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,
im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,
re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24,re_X2_0,im_X2_0,re_X2_1,im_X2_1,re_X2_2,im_X2_2,re_X2_3,im_X2_3,re_X2_4,im_X2_4,
re_X2_5,im_X2_5,re_X2_6,im_X2_6,re_X2_7,im_X2_7,re_X2_8,im_X2_8,re_X2_9,im_X2_9,re_X2_10,im_X2_10,re_X2_11,im_X2_11,re_X2_12,im_X2_12,re_X2_13,im_X2_13,re_X2_14,im_X2_14,re_X2_15,im_X2_15,
re_X2_16,im_X2_16,re_X2_17,im_X2_17,re_X2_18,im_X2_18,re_X2_19,im_X2_19,re_X2_20,im_X2_20,re_X2_21,im_X2_21,re_X2_22,im_X2_22,re_X2_23,im_X2_23,re_X2_24,im_X2_24,re_X_0,im_X_0,re_X_1,im_X_1,re_X_2,im_X_2,re_X_3,im_X_3,re_X_4,im_X_4,re_X_5,im_X_5,re_X_6,im_X_6,re_X_7,im_X_7,re_X_8,im_X_8,re_X_9,im_X_9,re_X_10,im_X_10,
re_X_11,im_X_11,re_X_12,im_X_12,re_X_13,im_X_13,re_X_14,im_X_14,re_X_15,im_X_15,re_X_16,im_X_16,re_X_17,im_X_17,re_X_18,im_X_18,re_X_19,im_X_19,re_X_20,im_X_20,re_X_21,im_X_21,
re_X_22,im_X_22,re_X_23,im_X_23,re_X_24,im_X_24,re_X_25,im_X_25,re_X_26,im_X_26,re_X_27,im_X_27,re_X_28,im_X_28,re_X_29,im_X_29,re_X_30,im_X_30,re_X_31,im_X_31,re_X_32,im_X_32,
re_X_33,im_X_33,re_X_34,im_X_34,re_X_35,im_X_35,re_X_36,im_X_36,re_X_37,im_X_37,re_X_38,im_X_38,re_X_39,im_X_39,re_X_40,im_X_40,re_X_41,im_X_41,re_X_42,im_X_42,re_X_43,im_X_43,
re_X_44,im_X_44,re_X_45,im_X_45,re_X_46,im_X_46,re_X_47,im_X_47,re_X_48,im_X_48,re_X_49,im_X_49);


input signed [16:0] re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,
im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,
re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24,re_X2_0,im_X2_0,re_X2_1,im_X2_1,re_X2_2,im_X2_2,re_X2_3,im_X2_3,re_X2_4,im_X2_4,
re_X2_5,im_X2_5,re_X2_6,im_X2_6,re_X2_7,im_X2_7,re_X2_8,im_X2_8,re_X2_9,im_X2_9,re_X2_10,im_X2_10,re_X2_11,im_X2_11,re_X2_12,im_X2_12,re_X2_13,im_X2_13,re_X2_14,im_X2_14,re_X2_15,im_X2_15,
re_X2_16,im_X2_16,re_X2_17,im_X2_17,re_X2_18,im_X2_18,re_X2_19,im_X2_19,re_X2_20,im_X2_20,re_X2_21,im_X2_21,re_X2_22,im_X2_22,re_X2_23,im_X2_23,re_X2_24,im_X2_24;

output reg signed [15:0] re_X_0,im_X_0,re_X_1,im_X_1,re_X_2,im_X_2,re_X_3,im_X_3,re_X_4,im_X_4,re_X_5,im_X_5,re_X_6,im_X_6,re_X_7,im_X_7,re_X_8,im_X_8,re_X_9,im_X_9,re_X_10,im_X_10,
re_X_11,im_X_11,re_X_12,im_X_12,re_X_13,im_X_13,re_X_14,im_X_14,re_X_15,im_X_15,re_X_16,im_X_16,re_X_17,im_X_17,re_X_18,im_X_18,re_X_19,im_X_19,re_X_20,im_X_20,re_X_21,im_X_21,
re_X_22,im_X_22,re_X_23,im_X_23,re_X_24,im_X_24,re_X_25,im_X_25,re_X_26,im_X_26,re_X_27,im_X_27,re_X_28,im_X_28,re_X_29,im_X_29,re_X_30,im_X_30,re_X_31,im_X_31,re_X_32,im_X_32,
re_X_33,im_X_33,re_X_34,im_X_34,re_X_35,im_X_35,re_X_36,im_X_36,re_X_37,im_X_37,re_X_38,im_X_38,re_X_39,im_X_39,re_X_40,im_X_40,re_X_41,im_X_41,re_X_42,im_X_42,re_X_43,im_X_43,
re_X_44,im_X_44,re_X_45,im_X_45,re_X_46,im_X_46,re_X_47,im_X_47,re_X_48,im_X_48,re_X_49,im_X_49;

input clk;

reg signed [31:0] m [295:0] ;
reg signed [14:0] n [295:0] ;
reg signed [18:0] p [99:0]  ;

wire signed [14:0] cos_0 , cos_7_2 , sin_7_2 , cos_14_4 , sin_14_4 , cos_21_6 , sin_21_6 , cos_28_8 , sin_28_8 , cos_36 , sin_36 , cos_43_2 , sin_43_2 , cos_50_4 , sin_50_4 , cos_57_2 , sin_57_2 
, cos_64_8 , sin_64_8 , cos_72 , sin_72 , cos_79_2 , sin_79_2 , cos_86_4 , sin_86_4 , cos_93_6 , sin_93_6 , cos_100_8 , sin_100_8 , cos_108 , sin_108 , cos_115_2 , sin_115_2 , cos_122_4 , sin_122_4,
cos_129_6 , sin_129_6 , cos_136_8 , sin_136_8 , cos_144 , sin_144 , cos_151_2 ,sin_151_2 , cos_158_4 , sin_158_4 , cos_165_6 , sin_165_6 , cos_172_8 , sin_172_8 ,cos_187_2,sin_187_2,cos_194_4,sin_194_4,
cos_201_6,sin_201_6,cos_208_8,sin_208_8,cos_216,sin_216,cos_223_2,sin_223_2,cos_230_4,sin_230_4,cos_237_6,sin_237_6,cos_244_8,sin_244_8,cos_252,sin_252,cos_259_2,sin_259_2,cos_266_4,sin_266_4,cos_273_6,
sin_273_6,cos_280_8,sin_280_8,cos_288,sin_288,cos_295_2,sin_295_2,cos_302_4,sin_302_4,cos_309_6,sin_309_6,cos_316_8,sin_316_8,cos_324,sin_324,cos_331_2,sin_331_2,cos_338_4,sin_338_4,cos_345_6,sin_345_6,cos_352_8,sin_352_8;

wire signed [2:0] div_2 ;

assign cos_0     ='b011111111111111;
assign cos_7_2   ='b011111101111110;
assign sin_7_2   ='b000100000000101;
assign cos_14_4  ='b011110111111101;
assign sin_14_4  ='b000111111101010;
assign cos_21_6  ='b011101110000001;
assign sin_21_6  ='b001011110001111;
assign cos_28_8  ='b011100000010101;
assign sin_28_8  ='b001111011010101;
assign cos_36    ='b011001111000110;
assign sin_36    ='b010010110011110;
assign cos_43_2  ='b010111010100111;
assign sin_43_2  ='b010101111001111;
assign cos_50_4  ='b010100011001011;
assign sin_50_4  ='b011000101010000;
assign cos_57_6  ='b010001001001010;
assign sin_57_6  ='b011011000001001;
assign cos_64_8  ='b001101100111111;
assign sin_64_8  ='b011100111101000;
assign cos_72    ='b001001111000110;
assign sin_72    ='b011110011011110;
assign cos_79_2  ='b000101111111110;
assign sin_79_2  ='b011111011011101;
assign cos_86_4  ='b000010000000100;
assign sin_86_4  ='b011111111011111;
assign cos_93_6  ='b111101111111100;
assign sin_93_6  ='b011111111011111;
assign cos_100_8 ='b111010000000100;
assign sin_100_8 ='b011111011011100;
assign cos_108   ='b110110000111010;
assign sin_108   ='b011110011011110;
assign cos_115_2 ='b110010011000010;
assign sin_115_2 ='b011100111101000;
assign cos_122_4 ='b101110110110110;
assign sin_122_4 ='b011011000001001;
assign cos_129_6 ='b101011100110101;
assign sin_129_6 ='b011000101001111;
assign cos_136_8 ='b101000101011001;
assign sin_136_8 ='b010101111001111;
assign cos_144   ='b100110000111010;
assign sin_144   ='b010010110011110;
assign cos_151_2 ='b100011111101011;
assign sin_151_2 ='b001111011010101;
assign cos_158_4 ='b100010010000000;
assign sin_158_4 ='b001011110001110;
assign cos_165_6 ='b100001000000011;
assign sin_165_6 ='b000111111101010;
assign cos_172_8 ='b100000010000010;
assign sin_172_8 ='b000100000000101;
assign cos_187_2 ='b100000010000010;
assign sin_187_2 ='b111011111111011;
assign cos_194_4 ='b100001000000011;
assign sin_194_4 ='b111000000010110;
assign cos_201_6 ='b100010010000000;
assign sin_201_6 ='b110100001110010;
assign cos_208_8 ='b100011111101011;
assign sin_208_8 ='b110000100101011;
assign cos_216   ='b100110000111010;
assign sin_216   ='b101101001100010;
assign cos_223_2 ='b101000101011001;
assign sin_223_2 ='b101010000110001;
assign cos_230_4 ='b101011100110101;
assign sin_230_4 ='b100111010110001;
assign cos_237_6 ='b101110110110110;
assign sin_237_6 ='b100100111110111;
assign cos_244_8 ='b110010011000010;
assign sin_244_8 ='b100011000011000;
assign cos_252   ='b110110000111010;
assign sin_252   ='b100001100100010;
assign cos_259_2 ='b111010000000100;
assign sin_259_2 ='b100000100100100;
assign cos_266_4 ='b111101111111100;
assign sin_266_4 ='b100000000100001;
assign cos_273_6 ='b000010000000100;
assign sin_273_6 ='b100000000100001;
assign cos_280_8 ='b000101111111110;
assign sin_280_8 ='b100000100100011;
assign cos_288   ='b001001111000110;
assign sin_288   ='b100001100100010;
assign cos_295_2 ='b001101100111111;
assign sin_295_2 ='b100011000011000;
assign cos_302_4 ='b010001001001010;
assign sin_302_4 ='b100100111110111;
assign cos_309_6 ='b010100011001011;
assign sin_309_6 ='b100111010110000;
assign cos_316_8 ='b010111010100111;
assign sin_316_8 ='b101010000110001;
assign cos_324   ='b011001111000110;
assign sin_324   ='b101101001100010;
assign cos_331_2 ='b011100000010101;
assign sin_331_2 ='b110000100101011;
assign cos_338_4 ='b011101110000001;
assign sin_338_4 ='b110100001110001;
assign cos_345_6 ='b011110111111101;
assign sin_345_6 ='b111000000010110;
assign cos_352_8 ='b011111101111110;
assign sin_352_8 ='b111011111111011;
assign div_2     ='b010;


always@(posedge clk)
begin

/////////////////////////////////////////////////////////////////// output of re_X_0

m[0]= (re_X1_0 * cos_0);
m[1]= (re_X2_0 * cos_0);

n[0]= m[0][31:17] + m[0][16];
n[1]= m[1][31:17] + m[1][16];

////////////////////////////////////////////////////////////////// output of im_X_0

m[2]= (im_X1_0 * cos_0);
m[3]= (im_X2_0 * cos_0); 

n[2]= m[2][31:17] + m[2][16];
n[3]= m[3][31:17] + m[3][16];

///////////////////////////////////////////////////////////////// output of re_X_1

m[4]= (re_X1_1 * cos_0);
m[5]= (re_X2_1 * cos_7_2);
m[6]= (im_X2_1 * sin_7_2);

n[4]= m[4][31:17] + m[4][16];
n[5]= m[5][31:17] + m[5][16];
n[6]= m[6][31:17] + m[6][16];

///////////////////////////////////////////////////////////////// output of im_X_1

m[7]= (im_X1_1 * cos_0);
m[8]= (im_X2_1 * cos_7_2);
m[9]= (re_X2_1 * sin_7_2);

n[7]= m[7][31:17] + m[7][16];
n[8]= m[8][31:17] + m[8][16];
n[9]= m[9][31:17] + m[9][16];

/////////////////////////////////////////////////////////////////output of re_X_2

m[10]= (re_X1_2 * cos_0);
m[11]= (re_X2_2 * cos_14_4);
m[12]= (im_X2_2 * sin_14_4);

n[10]= m[10][31:17] + m[10][16];
n[11]= m[11][31:17] + m[11][16];
n[12]= m[12][31:17] + m[12][16];

////////////////////////////////////////////////////////////////output of im_X_2

m[13]= (im_X1_2 * cos_0);
m[14]= (im_X2_2 * cos_14_4);
m[15]= (re_X2_2 * sin_14_4);

n[13]= m[13][31:17] + m[13][16];
n[14]= m[14][31:17] + m[14][16];
n[15]= m[15][31:17] + m[15][16];

////////////////////////////////////////////////////////////////output of re_X_3

m[16]= (re_X1_3 * cos_0);
m[17]= (re_X2_3 * cos_21_6);
m[18]= (im_X2_3 * sin_21_6);

n[16]= m[16][31:17] + m[16][16];
n[17]= m[17][31:17] + m[17][16];
n[18]= m[18][31:17] + m[18][16];

////////////////////////////////////////////////////////////////output of im_X_3

m[19]= (im_X1_3 * cos_0);
m[20]= (im_X2_3 * cos_21_6);
m[21]= (re_X2_3 * sin_21_6);

n[19]= m[19][31:17] + m[19][16];
n[20]= m[20][31:17] + m[20][16];
n[21]= m[21][31:17] + m[21][16];

//////////////////////////////////////////////////////////////////output of re_X_4

m[22]= (re_X1_4 * cos_0);
m[23]= (re_X2_4 * cos_28_8);
m[24]= (im_X2_4 * sin_28_8);

n[22]= m[22][31:17] + m[22][16];
n[23]= m[23][31:17] + m[23][16];
n[24]= m[24][31:17] + m[24][16];

/////////////////////////////////////////////////////////////////output of im_X_4

m[25]= (im_X1_4 * cos_0);
m[26]= (im_X2_4 * cos_28_8);
m[27]= (re_X2_4 * sin_28_8);

n[25]= m[25][31:17] + m[25][16];
n[26]= m[26][31:17] + m[26][16];
n[27]= m[27][31:17] + m[27][16];

/////////////////////////////////////////////////////////////////output of re_X_5

m[28]= (re_X1_5 * cos_0);
m[29]= (re_X2_5 * cos_36);
m[30]= (im_X2_5 * sin_36);

n[28]= m[28][31:17] + m[28][16];
n[29]= m[29][31:17] + m[29][16];
n[30]= m[30][31:17] + m[30][16];

//////////////////////////////////////////////////////////////////output of im_X_5

m[31]= (im_X1_5 * cos_0);
m[32]= (im_X2_5 * cos_36);
m[33]= (re_X2_5 * sin_36);

n[31]= m[31][31:17] + m[31][16];
n[32]= m[32][31:17] + m[32][16];
n[33]= m[33][31:17] + m[33][16];

////////////////////////////////////////////////////////////////output of re_X_6

m[34]= (re_X1_6 * cos_0);
m[35]= (re_X2_6 * cos_43_2);
m[36]= (im_X2_6 * sin_43_2);

n[34]= m[34][31:17] + m[34][16];
n[35]= m[35][31:17] + m[35][16];
n[36]= m[36][31:17] + m[36][16];

///////////////////////////////////////////////////////////////output of im_X_6

m[37]= (im_X1_6 * cos_0);
m[38]= (im_X2_6 * cos_43_2);
m[39]= (re_X2_6 * sin_43_2);

n[37]= m[37][31:17] + m[37][16];
n[38]= m[38][31:17] + m[38][16];
n[39]= m[39][31:17] + m[39][16];

///////////////////////////////////////////////////////////////output of re_X_7

m[40]= (re_X1_7 * cos_0);
m[41]= (re_X2_7 * cos_50_4);
m[42]= (im_X2_7 * sin_50_4);

n[40]= m[40][31:17] + m[40][16];
n[41]= m[41][31:17] + m[41][16];
n[42]= m[42][31:17] + m[42][16];

///////////////////////////////////////////////////////////////output of im_X_7

m[43]= (im_X1_7 * cos_0);
m[44]= (im_X2_7 * cos_50_4);
m[45]= (re_X2_7 * sin_50_4);

n[43]= m[43][31:17] + m[43][16];
n[44]= m[44][31:17] + m[44][16];
n[45]= m[45][31:17] + m[45][16];

///////////////////////////////////////////////////////////////output of re_X_8

m[46]= (re_X1_8 * cos_0);
m[47]= (re_X2_8 * cos_57_6);
m[48]= (im_X2_8 * sin_57_6);

n[46]= m[46][31:17] + m[46][16];
n[47]= m[47][31:17] + m[47][16];
n[48]= m[48][31:17] + m[48][16];

///////////////////////////////////////////////////////////////output of im_X_8

m[49]= (im_X1_8 * cos_0);
m[50]= (im_X2_8 * cos_57_6);
m[51]= (re_X2_8 * sin_57_6);

n[49]= m[49][31:17] + m[49][16];
n[50]= m[50][31:17] + m[50][16];
n[51]= m[51][31:17] + m[51][16];

///////////////////////////////////////////////////////////////output of re_X_9

m[52]= (re_X1_9 * cos_0);
m[53]= (re_X2_9 * cos_64_8);
m[54]= (im_X2_9 * sin_64_8);

n[52]= m[52][31:17] + m[52][16];
n[53]= m[53][31:17] + m[53][16];
n[54]= m[54][31:17] + m[54][16];

///////////////////////////////////////////////////////////////output of im_X_9

m[55]= (im_X1_9 * cos_0);
m[56]= (im_X2_9 * cos_64_8);
m[57]= (re_X2_9 * sin_64_8);

n[55]= m[55][31:17] + m[55][16];
n[56]= m[56][31:17] + m[56][16];
n[57]= m[57][31:17] + m[57][16];

///////////////////////////////////////////////////////////////output of re_X_10

m[58]= (re_X1_10 * cos_0);
m[59]= (re_X2_10 * cos_72);
m[60]= (im_X2_10 * sin_72);

n[58]= m[58][31:17] + m[58][16];
n[59]= m[59][31:17] + m[59][16];
n[60]= m[60][31:17] + m[60][16];

///////////////////////////////////////////////////////////////output of im_X_10

m[61]= (im_X1_10 * cos_0);
m[62]= (im_X2_10 * cos_72);
m[63]= (re_X2_10 * sin_72);

n[61]= m[61][31:17] + m[61][16];
n[62]= m[62][31:17] + m[62][16];
n[63]= m[63][31:17] + m[63][16];

///////////////////////////////////////////////////////////////output of re_X_11

m[64]= (re_X1_11 * cos_0);
m[65]= (re_X2_11 * cos_79_2);
m[66]= (im_X2_11 * sin_79_2);

n[64]= m[64][31:17] + m[64][16];
n[65]= m[65][31:17] + m[65][16];
n[66]= m[66][31:17] + m[66][16];

///////////////////////////////////////////////////////////////output of im_X_11

m[67]= (im_X1_11 * cos_0);
m[68]= (im_X2_11 * cos_79_2);
m[69]= (re_X2_11 * sin_79_2);

n[67]= m[67][31:17] + m[67][16];
n[68]= m[68][31:17] + m[68][16];
n[69]= m[69][31:17] + m[69][16];

///////////////////////////////////////////////////////////////output of re_X_12

m[70]= (re_X1_12 * cos_0);
m[71]= (re_X2_12 * cos_86_4);
m[72]= (im_X2_12 * sin_86_4);

n[70]= m[70][31:17] + m[70][16];
n[71]= m[71][31:17] + m[71][16];
n[72]= m[72][31:17] + m[72][16];

///////////////////////////////////////////////////////////////output of im_X_12

m[73]= (im_X1_12 * cos_0);
m[74]= (im_X2_12 * cos_86_4);
m[75]= (re_X2_12 * sin_86_4);

n[73]= m[73][31:17] + m[73][16];
n[74]= m[74][31:17] + m[74][16];
n[75]= m[75][31:17] + m[75][16];

///////////////////////////////////////////////////////////////output of re_X_13

m[76]= (re_X1_13 * cos_0);
m[77]= (re_X2_13 * cos_93_6);
m[78]= (im_X2_13 * sin_93_6);

n[76]= m[76][31:17] + m[76][16];
n[77]= m[77][31:17] + m[77][16];
n[78]= m[78][31:17] + m[78][16];

///////////////////////////////////////////////////////////////output of im_X_13

m[79]= (im_X1_13 * cos_0);
m[80]= (im_X2_13 * cos_93_6);
m[81]= (re_X2_13 * sin_93_6);

n[79]= m[79][31:17] + m[79][16];
n[80]= m[80][31:17] + m[80][16];
n[81]= m[81][31:17] + m[81][16];

///////////////////////////////////////////////////////////////output of re_X_14

m[82]= (re_X1_14 * cos_0);
m[83]= (re_X2_14 * cos_100_8);
m[84]= (im_X2_14 * sin_100_8);

n[82]= m[82][31:17] + m[82][16];
n[83]= m[83][31:17] + m[83][16];
n[84]= m[84][31:17] + m[84][16];

///////////////////////////////////////////////////////////////output of im_X_14

m[85]= (im_X1_14 * cos_0);
m[86]= (im_X2_14 * cos_100_8);
m[87]= (re_X2_14 * sin_100_8);

n[85]= m[85][31:17] + m[85][16];
n[86]= m[86][31:17] + m[86][16];
n[87]= m[87][31:17] + m[87][16];


///////////////////////////////////////////////////////////////output of re_X_15

m[88]= (re_X1_15 * cos_0);
m[89]= (re_X2_15 * cos_108);
m[90]= (im_X2_15 * sin_108);

n[88]= m[88][31:17] + m[88][16];
n[89]= m[89][31:17] + m[89][16];
n[90]= m[90][31:17] + m[90][16];

///////////////////////////////////////////////////////////////output of im_X_15

m[91]= (im_X1_15 * cos_0);
m[92]= (im_X2_15 * cos_108);
m[93]= (re_X2_15 * sin_108);

n[91]= m[91][31:17] + m[91][16];
n[92]= m[92][31:17] + m[92][16];
n[93]= m[93][31:17] + m[93][16];


///////////////////////////////////////////////////////////////output of re_X_16

m[94]= (re_X1_16 * cos_0);
m[95]= (re_X2_16 * cos_115_2);
m[96]= (im_X2_16 * sin_115_2);

n[94]= m[94][31:17] + m[94][16];
n[95]= m[95][31:17] + m[95][16];
n[96]= m[96][31:17] + m[96][16];

///////////////////////////////////////////////////////////////output of im_X_16

m[97]= (im_X1_16 * cos_0);
m[98]= (im_X2_16 * cos_115_2);
m[99]= (re_X2_16 * sin_115_2);

n[97]= m[97][31:17] + m[97][16];
n[98]= m[98][31:17] + m[98][16];
n[99]= m[99][31:17] + m[99][16];

///////////////////////////////////////////////////////////////output of re_X_17

m[100]= (re_X1_17 * cos_0);
m[101]= (re_X2_17 * cos_122_4);
m[102]= (im_X2_17 * sin_122_4);

n[100]= m[100][31:17] + m[100][16];
n[101]= m[101][31:17] + m[101][16];
n[102]= m[102][31:17] + m[102][16];

///////////////////////////////////////////////////////////////output of im_X_17

m[103]= (im_X1_17 * cos_0);
m[104]= (im_X2_17 * cos_122_4);
m[105]= (re_X2_17 * sin_122_4);

n[103]= m[103][31:17] + m[103][16];
n[104]= m[104][31:17] + m[104][16];
n[105]= m[105][31:17] + m[105][16];

///////////////////////////////////////////////////////////////output of re_X_18

m[106]= (re_X1_18 * cos_0);
m[107]= (re_X2_18 * cos_129_6);
m[108]= (im_X2_18 * sin_129_6);

n[106]= m[106][31:17] + m[106][16];
n[107]= m[107][31:17] + m[107][16];
n[108]= m[108][31:17] + m[108][16];

///////////////////////////////////////////////////////////////output of im_X_18

m[109]= (im_X1_18 * cos_0);
m[110]= (im_X2_18 * cos_129_6);
m[111]= (re_X2_18 * sin_129_6);

n[109]= m[109][31:17] + m[109][16];
n[110]= m[110][31:17] + m[110][16];
n[111]= m[111][31:17] + m[111][16];

///////////////////////////////////////////////////////////////output of re_X_19

m[112]= (re_X1_19 * cos_0);
m[113]= (re_X2_19 * cos_136_8);
m[114]= (im_X2_19 * sin_136_8);

n[112]= m[112][31:17] + m[112][16];
n[113]= m[113][31:17] + m[113][16];
n[114]= m[114][31:17] + m[114][16];

///////////////////////////////////////////////////////////////output of im_X_19

m[115]= (im_X1_19 * cos_0);
m[116]= (im_X2_19 * cos_136_8);
m[117]= (re_X2_19 * sin_136_8);

n[115]= m[115][31:17] + m[115][16];
n[116]= m[116][31:17] + m[116][16];
n[117]= m[117][31:17] + m[117][16];

///////////////////////////////////////////////////////////////output of re_X_20

m[118]= (re_X1_20 * cos_0);
m[119]= (re_X2_20 * cos_144);
m[120]= (im_X2_20 * sin_144);

n[118]= m[118][31:17] + m[118][16];
n[119]= m[119][31:17] + m[119][16];
n[120]= m[120][31:17] + m[120][16];

///////////////////////////////////////////////////////////////output of im_X_20

m[121]= (im_X1_20 * cos_0);
m[122]= (im_X2_20 * cos_144);
m[123]= (re_X2_20 * sin_144);

n[121]= m[121][31:17] + m[121][16];
n[122]= m[122][31:17] + m[122][16];
n[123]= m[123][31:17] + m[123][16];

///////////////////////////////////////////////////////////////output of re_X_21

m[124]= (re_X1_21 * cos_0);
m[125]= (re_X2_21 * cos_151_2);
m[126]= (im_X2_21 * sin_151_2);

n[124]= m[124][31:17] + m[124][16];
n[125]= m[125][31:17] + m[125][16];
n[126]= m[126][31:17] + m[126][16];

///////////////////////////////////////////////////////////////output of im_X_21

m[127]= (im_X1_21 * cos_0);
m[128]= (im_X2_21 * cos_151_2);
m[129]= (re_X2_21 * sin_151_2);

n[127]= m[127][31:17] + m[127][16];
n[128]= m[128][31:17] + m[128][16];
n[129]= m[129][31:17] + m[129][16];

///////////////////////////////////////////////////////////////output of re_X_22

m[130]= (re_X1_22 * cos_0);
m[131]= (re_X2_22 * cos_158_4);
m[132]= (im_X2_22 * sin_158_4);

n[130]= m[130][31:17] + m[130][16];
n[131]= m[131][31:17] + m[131][16];
n[132]= m[132][31:17] + m[132][16];

///////////////////////////////////////////////////////////////output of im_X_22

m[133]= (im_X1_22 * cos_0);
m[134]= (im_X2_22 * cos_158_4);
m[135]= (re_X2_22 * sin_158_4);

n[133]= m[133][31:17] + m[133][16];
n[134]= m[134][31:17] + m[134][16];
n[135]= m[135][31:17] + m[135][16];

///////////////////////////////////////////////////////////////output of re_X_23

m[136]= (re_X1_23 * cos_0);
m[137]= (re_X2_23 * cos_165_6);
m[138]= (im_X2_23 * sin_165_6);

n[136]= m[136][31:17] + m[136][16];
n[137]= m[137][31:17] + m[137][16];
n[138]= m[138][31:17] + m[138][16];

///////////////////////////////////////////////////////////////output of im_X_23

m[139]= (im_X1_23 * cos_0);
m[140]= (im_X2_23 * cos_165_6);
m[141]= (re_X2_23 * sin_165_6);

n[139]= m[139][31:17] + m[139][16];
n[140]= m[140][31:17] + m[140][16];
n[141]= m[141][31:17] + m[141][16];

///////////////////////////////////////////////////////////////output of re_X_24

m[142]= (re_X1_24 * cos_0);
m[143]= (re_X2_24 * cos_172_8);
m[144]= (im_X2_24 * sin_172_8);

n[142]= m[142][31:17] + m[142][16];
n[143]= m[143][31:17] + m[143][16];
n[144]= m[144][31:17] + m[144][16];

///////////////////////////////////////////////////////////////output of im_X_24

m[145]= (im_X1_24 * cos_0);
m[146]= (im_X2_24 * cos_172_8);
m[147]= (re_X2_24 * sin_172_8);

n[145]= m[145][31:17] + m[145][16];
n[146]= m[146][31:17] + m[146][16];
n[147]= m[147][31:17] + m[147][16];

///////////////////////////////////////////////////////////////output of re_X_25

m[148]= (re_X1_0 * cos_0);
m[149]= (re_X2_0 * cos_0);

n[148]= m[148][31:17] + m[148][16];
n[149]= m[149][31:17] + m[149][16];

///////////////////////////////////////////////////////////////output of im_X_25

m[150]= (im_X1_0 * cos_0);
m[151]= (im_X2_0 * cos_0); 

n[150]= m[150][31:17] + m[150][16];
n[151]= m[151][31:17] + m[151][16];

//////////////////////////////////////////////////////////////// output of re_X_26

m[152]= (re_X1_1 * cos_0);
m[153]= (re_X2_1 * cos_187_2);
m[154]= (im_X2_1 * sin_187_2);

n[152]= m[152][31:17] + m[152][16];
n[153]= m[153][31:17] + m[153][16];
n[154]= m[154][31:17] + m[154][16];

///////////////////////////////////////////////////////////////// output of im_X_26

m[155]= (im_X1_1 * cos_0);
m[156]= (im_X2_1 * cos_187_2);
m[157]= (re_X2_1 * sin_187_2);

n[155]= m[155][31:17] + m[155][16];
n[156]= m[156][31:17] + m[156][16];
n[157]= m[157][31:17] + m[157][16];

///////////////////////////////////////////////////////////////// output of re_X_27

m[158]= (re_X1_2 * cos_0);
m[159]= (re_X2_2 * cos_194_4);
m[160]= (im_X2_2 * sin_194_4);

n[158]= m[158][31:17] + m[158][16];
n[159]= m[159][31:17] + m[159][16];
n[160]= m[160][31:17] + m[160][16];

///////////////////////////////////////////////////////////////// output of im_X_27

m[161]= (im_X1_2 * cos_0);
m[162]= (im_X2_2 * cos_194_4);
m[163]= (re_X2_2 * sin_194_4);

n[161]= m[161][31:17] + m[161][16];
n[162]= m[162][31:17] + m[162][16];
n[163]= m[163][31:17] + m[163][16];

///////////////////////////////////////////////////////////////// output of re_X_28

m[164]= (re_X1_3 * cos_0);
m[165]= (re_X2_3 * cos_201_6);
m[166]= (im_X2_3 * sin_201_6);

n[164]= m[164][31:17] + m[164][16];
n[165]= m[165][31:17] + m[165][16];
n[166]= m[166][31:17] + m[166][16];

///////////////////////////////////////////////////////////////// output of im_X_28

m[167]= (im_X1_3 * cos_0);
m[168]= (im_X2_3 * cos_201_6);
m[169]= (re_X2_3 * sin_201_6);

n[167]= m[167][31:17] + m[167][16];
n[168]= m[168][31:17] + m[168][16];
n[169]= m[169][31:17] + m[169][16];


///////////////////////////////////////////////////////////////// output of re_X_29

m[170]= (re_X1_4 * cos_0);
m[171]= (re_X2_4 * cos_208_8);
m[172]= (im_X2_4 * sin_208_8);

n[170]= m[170][31:17] + m[170][16];
n[171]= m[171][31:17] + m[171][16];
n[172]= m[172][31:17] + m[172][16];

///////////////////////////////////////////////////////////////// output of im_X_29

m[173]= (im_X1_4 * cos_0);
m[174]= (im_X2_4 * cos_208_8);
m[175]= (re_X2_4 * sin_208_8);

n[173]= m[173][31:17] + m[173][16];
n[174]= m[174][31:17] + m[174][16];
n[175]= m[175][31:17] + m[175][16];



///////////////////////////////////////////////////////////////// output of re_X_30

m[176]= (re_X1_5 * cos_0);
m[177]= (re_X2_5 * cos_216);
m[178]= (im_X2_5 * sin_216);

n[176]= m[176][31:17] + m[176][16];
n[177]= m[177][31:17] + m[177][16];
n[178]= m[178][31:17] + m[178][16];

///////////////////////////////////////////////////////////////// output of im_X_30

m[179]= (im_X1_5 * cos_0);
m[180]= (im_X2_5 * cos_216);
m[181]= (re_X2_5 * sin_216);

n[179]= m[179][31:17] + m[179][16];
n[180]= m[180][31:17] + m[180][16];
n[181]= m[181][31:17] + m[181][16];



///////////////////////////////////////////////////////////////// output of re_X_31

m[182]= (re_X1_6 * cos_0);
m[183]= (re_X2_6 * cos_223_2);
m[184]= (im_X2_6 * sin_223_2);

n[182]= m[182][31:17] + m[182][16];
n[183]= m[183][31:17] + m[183][16];
n[184]= m[184][31:17] + m[184][16];

///////////////////////////////////////////////////////////////// output of im_X_31

m[185]= (im_X1_6 * cos_0);
m[186]= (im_X2_6 * cos_223_2);
m[187]= (re_X2_6 * sin_223_2);

n[185]= m[185][31:17] + m[185][16];
n[186]= m[186][31:17] + m[186][16];
n[187]= m[187][31:17] + m[187][16];


///////////////////////////////////////////////////////////////// output of re_X_32

m[188]= (re_X1_7 * cos_0);
m[189]= (re_X2_7 * cos_230_4);
m[190]= (im_X2_7 * sin_230_4);

n[188]= m[188][31:17] + m[188][16];
n[189]= m[189][31:17] + m[189][16];
n[190]= m[190][31:17] + m[190][16];

///////////////////////////////////////////////////////////////// output of im_X_32

m[191]= (im_X1_7 * cos_0);
m[192]= (im_X2_7 * cos_230_4);
m[193]= (re_X2_7 * sin_230_4);

n[191]= m[191][31:17] + m[191][16];
n[192]= m[192][31:17] + m[192][16];
n[193]= m[193][31:17] + m[193][16];




///////////////////////////////////////////////////////////////// output of re_X_33

m[194]= (re_X1_8 * cos_0);
m[195]= (re_X2_8 * cos_237_6);
m[196]= (im_X2_8 * sin_237_6);

n[194]= m[194][31:17] + m[194][16];
n[195]= m[195][31:17] + m[195][16];
n[196]= m[196][31:17] + m[196][16];

///////////////////////////////////////////////////////////////// output of im_X_33

m[197]= (im_X1_8 * cos_0);
m[198]= (im_X2_8 * cos_237_6);
m[199]= (re_X2_8 * sin_237_6);

n[197]= m[197][31:17] + m[197][16];
n[198]= m[198][31:17] + m[198][16];
n[199]= m[199][31:17] + m[199][16];



///////////////////////////////////////////////////////////////// output of re_X_34

m[200]= (re_X1_9 * cos_0);
m[201]= (re_X2_9 * cos_244_8);
m[202]= (im_X2_9 * sin_244_8);

n[200]= m[200][31:17] + m[200][16];
n[201]= m[201][31:17] + m[201][16];
n[202]= m[202][31:17] + m[202][16];

///////////////////////////////////////////////////////////////// output of im_X_34

m[203]= (im_X1_9 * cos_0);
m[204]= (im_X2_9 * cos_244_8);
m[205]= (re_X2_9 * sin_244_8);

n[203]= m[203][31:17] + m[203][16];
n[204]= m[204][31:17] + m[204][16];
n[205]= m[205][31:17] + m[205][16];

///////////////////////////////////////////////////////////////// output of re_X_35

m[206]= (re_X1_10 * cos_0);
m[207]= (re_X2_10 * cos_252);
m[208]= (im_X2_10 * sin_252);

n[206]= m[206][31:17] + m[206][16];
n[207]= m[207][31:17] + m[207][16];
n[208]= m[208][31:17] + m[208][16];

///////////////////////////////////////////////////////////////// output of im_X_35

m[209]= (im_X1_10 * cos_0);
m[210]= (im_X2_10 * cos_252);
m[211]= (re_X2_10 * sin_252);

n[209]= m[209][31:17] + m[209][16];
n[210]= m[210][31:17] + m[210][16];
n[211]= m[211][31:17] + m[211][16];


///////////////////////////////////////////////////////////////// output of re_X_36

m[212]= (re_X1_11 * cos_0);
m[213]= (re_X2_11 * cos_259_2);
m[214]= (im_X2_11 * sin_259_2);

n[212]= m[212][31:17] + m[212][16];
n[213]= m[213][31:17] + m[213][16];
n[214]= m[214][31:17] + m[214][16];

///////////////////////////////////////////////////////////////// output of im_X_36

m[215]= (im_X1_11 * cos_0);
m[216]= (im_X2_11 * cos_259_2);
m[217]= (re_X2_11 * sin_259_2);

n[215]= m[215][31:17] + m[215][16];
n[216]= m[216][31:17] + m[216][16];
n[217]= m[217][31:17] + m[217][16];


///////////////////////////////////////////////////////////////// output of re_X_37

m[218]= (re_X1_12 * cos_0);
m[219]= (re_X2_12 * cos_266_4);
m[220]= (im_X2_12 * sin_266_4);

n[218]= m[218][31:17] + m[218][16];
n[219]= m[219][31:17] + m[219][16];
n[220]= m[220][31:17] + m[220][16];

///////////////////////////////////////////////////////////////// output of im_X_37

m[221]= (im_X1_12 * cos_0);
m[222]= (im_X2_12 * cos_266_4);
m[223]= (re_X2_12 * sin_266_4);

n[221]= m[221][31:17] + m[221][16];
n[222]= m[222][31:17] + m[222][16];
n[223]= m[223][31:17] + m[223][16];


///////////////////////////////////////////////////////////////// output of re_X_38

m[224]= (re_X1_13 * cos_0);
m[225]= (re_X2_13 * cos_273_6);
m[226]= (im_X2_13 * sin_273_6);

n[224]= m[224][31:17] + m[224][16];
n[225]= m[225][31:17] + m[225][16];
n[226]= m[226][31:17] + m[226][16];

///////////////////////////////////////////////////////////////// output of im_X_38

m[227]= (im_X1_13 * cos_0);
m[228]= (im_X2_13 * cos_273_6);
m[229]= (re_X2_13 * sin_273_6);

n[227]= m[227][31:17] + m[227][16];
n[228]= m[228][31:17] + m[228][16];
n[229]= m[229][31:17] + m[229][16];


///////////////////////////////////////////////////////////////// output of re_X_39

m[230]= (re_X1_14 * cos_0);
m[231]= (re_X2_14 * cos_280_8);
m[232]= (im_X2_14 * sin_280_8);

n[230]= m[230][31:17] + m[230][16];
n[231]= m[231][31:17] + m[231][16];
n[232]= m[232][31:17] + m[232][16];

///////////////////////////////////////////////////////////////// output of im_X_39

m[233]= (im_X1_14 * cos_0);
m[234]= (im_X2_14 * cos_280_8);
m[235]= (re_X2_14 * sin_280_8);

n[233]= m[233][31:17] + m[233][16];
n[234]= m[234][31:17] + m[234][16];
n[235]= m[235][31:17] + m[235][16];


///////////////////////////////////////////////////////////////// output of re_X_40

m[236]= (re_X1_15 * cos_0);
m[237]= (re_X2_15 * cos_288);
m[238]= (im_X2_15 * sin_288);

n[236]= m[236][31:17] + m[236][16];
n[237]= m[237][31:17] + m[237][16];
n[238]= m[238][31:17] + m[238][16];

///////////////////////////////////////////////////////////////// output of im_X_40

m[239]= (im_X1_15 * cos_0);
m[240]= (im_X2_15 * cos_288);
m[241]= (re_X2_15 * sin_288);

n[239]= m[239][31:17] + m[239][16];
n[240]= m[240][31:17] + m[240][16];
n[241]= m[241][31:17] + m[241][16];


///////////////////////////////////////////////////////////////// output of re_X_41

m[242]= (re_X1_16 * cos_0);
m[243]= (re_X2_16 * cos_295_2);
m[244]= (im_X2_16 * sin_295_2);

n[242]= m[242][31:17] + m[242][16];
n[243]= m[243][31:17] + m[243][16];
n[244]= m[244][31:17] + m[244][16];

///////////////////////////////////////////////////////////////// output of im_X_41

m[245]= (im_X1_16 * cos_0);
m[246]= (im_X2_16 * cos_295_2);
m[247]= (re_X2_16 * sin_295_2);

n[245]= m[245][31:17] + m[245][16];
n[246]= m[246][31:17] + m[246][16];
n[247]= m[247][31:17] + m[247][16];


///////////////////////////////////////////////////////////////// output of re_X_42

m[248]= (re_X1_17 * cos_0);
m[249]= (re_X2_17 * cos_302_4);
m[250]= (im_X2_17 * sin_302_4);

n[248]= m[248][31:17] + m[248][16];
n[249]= m[249][31:17] + m[249][16];
n[250]= m[250][31:17] + m[250][16];

///////////////////////////////////////////////////////////////// output of im_X_42

m[251]= (im_X1_17 * cos_0);
m[252]= (im_X2_17 * cos_302_4);
m[253]= (re_X2_17 * sin_302_4);

n[251]= m[251][31:17] + m[251][16];
n[252]= m[252][31:17] + m[252][16];
n[253]= m[253][31:17] + m[253][16];


///////////////////////////////////////////////////////////////// output of re_X_43

m[254]= (re_X1_18 * cos_0);
m[255]= (re_X2_18 * cos_309_6);
m[256]= (im_X2_18 * sin_309_6);

n[254]= m[254][31:17] + m[254][16];
n[255]= m[255][31:17] + m[255][16];
n[256]= m[256][31:17] + m[256][16];

///////////////////////////////////////////////////////////////// output of im_X_43

m[257]= (im_X1_18 * cos_0);
m[258]= (im_X2_18 * cos_309_6);
m[259]= (re_X2_18 * sin_309_6);

n[257]= m[257][31:17] + m[257][16];
n[258]= m[258][31:17] + m[258][16];
n[259]= m[259][31:17] + m[259][16];


///////////////////////////////////////////////////////////////// output of re_X_44

m[260]= (re_X1_19 * cos_0);
m[261]= (re_X2_19 * cos_316_8);
m[262]= (im_X2_19 * sin_316_8);

n[260]= m[260][31:17] + m[260][16];
n[261]= m[261][31:17] + m[261][16];
n[262]= m[262][31:17] + m[262][16];

///////////////////////////////////////////////////////////////// output of im_X_44

m[263]= (im_X1_19 * cos_0);
m[264]= (im_X2_19 * cos_316_8);
m[265]= (re_X2_19 * sin_316_8);

n[263]= m[263][31:17] + m[263][16];
n[264]= m[264][31:17] + m[264][16];
n[265]= m[265][31:17] + m[265][16];


///////////////////////////////////////////////////////////////// output of re_X_45

m[266]= (re_X1_20 * cos_0);
m[267]= (re_X2_20 * cos_324);
m[268]= (im_X2_20 * sin_324);

n[266]= m[266][31:17] + m[266][16];
n[267]= m[267][31:17] + m[267][16];
n[268]= m[268][31:17] + m[268][16];

///////////////////////////////////////////////////////////////// output of im_X_45

m[269]= (im_X1_20 * cos_0);
m[270]= (im_X2_20 * cos_324);
m[271]= (re_X2_20 * sin_324);

n[269]= m[269][31:17] + m[269][16];
n[270]= m[270][31:17] + m[270][16];
n[271]= m[271][31:17] + m[271][16];


///////////////////////////////////////////////////////////////// output of re_X_46

m[272]= (re_X1_21 * cos_0);
m[273]= (re_X2_21 * cos_331_2);
m[274]= (im_X2_21 * sin_331_2);

n[272]= m[272][31:17] + m[272][16];
n[273]= m[273][31:17] + m[273][16];
n[274]= m[274][31:17] + m[274][16];

///////////////////////////////////////////////////////////////// output of im_X_46

m[275]= (im_X1_21 * cos_0);
m[276]= (im_X2_21 * cos_331_2);
m[277]= (re_X2_21 * sin_331_2);

n[275]= m[275][31:17] + m[275][16];
n[276]= m[276][31:17] + m[276][16];
n[277]= m[277][31:17] + m[277][16];



///////////////////////////////////////////////////////////////// output of re_X_47

m[278]= (re_X1_22 * cos_0);
m[279]= (re_X2_22 * cos_338_4);
m[280]= (im_X2_22 * sin_338_4);

n[278]= m[278][31:17] + m[278][16];
n[279]= m[279][31:17] + m[279][16];
n[280]= m[280][31:17] + m[280][16];

///////////////////////////////////////////////////////////////// output of im_X_47

m[281]= (im_X1_22 * cos_0);
m[282]= (im_X2_22 * cos_338_4);
m[283]= (re_X2_22 * sin_338_4);

n[281]= m[281][31:17] + m[281][16];
n[282]= m[282][31:17] + m[282][16];
n[283]= m[283][31:17] + m[283][16];


///////////////////////////////////////////////////////////////// output of re_X_48

m[284]= (re_X1_23 * cos_0);
m[285]= (re_X2_23 * cos_345_6);
m[286]= (im_X2_23 * sin_345_6);

n[284]= m[284][31:17] + m[284][16];
n[285]= m[285][31:17] + m[285][16];
n[286]= m[286][31:17] + m[286][16];

///////////////////////////////////////////////////////////////// output of im_X_48

m[287]= (im_X1_23 * cos_0);
m[288]= (im_X2_23 * cos_345_6);
m[289]= (re_X2_23 * sin_345_6);

n[287]= m[287][31:17] + m[287][16];
n[288]= m[288][31:17] + m[288][16];
n[289]= m[289][31:17] + m[289][16];

///////////////////////////////////////////////////////////////// output of re_X_49

m[290]= (re_X1_24 * cos_0);
m[291]= (re_X2_24 * cos_352_8);
m[292]= (im_X2_24 * sin_352_8);

n[290]= m[290][31:17] + m[290][16];
n[291]= m[291][31:17] + m[291][16];
n[292]= m[292][31:17] + m[292][16];

///////////////////////////////////////////////////////////////// output of im_X_49

m[293]= (im_X1_24 * cos_0);
m[294]= (im_X2_24 * cos_352_8);
m[295]= (re_X2_24 * sin_352_8);

n[293]= m[293][31:17] + m[293][16];
n[294]= m[294][31:17] + m[294][16];
n[295]= m[295][31:17] + m[295][16];



//////////////////////////////////////////////////////////////////

p[0] = div_2*(n[0] + n[1]);
p[1] = div_2*(n[2] + n[3]);
p[2] = div_2*(n[4] + n[5] + n[6]);
p[3] = div_2*(n[7] + n[8] - n[9]);
p[4] = div_2*(n[10] + n[11] + n[12]);
p[5] = div_2*(n[13] + n[14] - n[15]);
p[6] = div_2*(n[16] + n[17] + n[18]);
p[7] = div_2*(n[19] + n[20] - n[21]);
p[8] = div_2*(n[22] + n[23] + n[24]);
p[9] = div_2*(n[25] + n[26] - n[27]);
p[10] = div_2*(n[28] + n[29] + n[30]);
p[11] = div_2*(n[31] + n[32] - n[33]);
p[12] = div_2*(n[34] + n[35] + n[36]);
p[13] = div_2*(n[37] + n[38] - n[39]);
p[14] = div_2*(n[40] + n[41] + n[42]);
p[15] = div_2*(n[43] + n[44] - n[45]);
p[16] = div_2*(n[46] + n[47] + n[48]);
p[17] = div_2*(n[49] + n[50] - n[51]);
p[18] = div_2*(n[52] + n[53] + n[54]);
p[19] = div_2*(n[55] + n[56] - n[57]);
p[20] = div_2*(n[58] + n[59] + n[60]);
p[21] = div_2*(n[61] + n[62] - n[63]);
p[22] = div_2*(n[64] + n[65] + n[66]);
p[23] = div_2*(n[67] + n[68] - n[69]);
p[24] = div_2*(n[70] + n[71] + n[72]);
p[25] = div_2*(n[73] + n[74] - n[75]);
p[26] = div_2*(n[76] + n[77] + n[78]);
p[27] = div_2*(n[79] + n[80] - n[81]);
p[28] = div_2*(n[82] + n[83] + n[84]);
p[29] = div_2*(n[85] + n[86] - n[87]);
p[30] = div_2*(n[88] + n[89] + n[90]);
p[31] = div_2*(n[91] + n[92] - n[93]);
p[32] = div_2*(n[94] + n[95] + n[96]);
p[33] = div_2*(n[97] + n[98] - n[99]);
p[34] = div_2*(n[100] + n[101] + n[102]);
p[35] = div_2*(n[103] + n[104] - n[105]);
p[36] = div_2*(n[106] + n[107] + n[108]);
p[37] = div_2*(n[109] + n[110] - n[111]);
p[38] = div_2*(n[112] + n[113] + n[114]);
p[39] = div_2*(n[115] + n[116] - n[117]);
p[40] = div_2*(n[118] + n[119] + n[120]);
p[41] = div_2*(n[121] + n[122] - n[123]);
p[42] = div_2*(n[124] + n[125] + n[126]);
p[43] = div_2*(n[127] + n[128] - n[129]);
p[44] = div_2*(n[130] + n[131] + n[132]);
p[45] = div_2*(n[133] + n[134] - n[135]);
p[46] = div_2*(n[136] + n[137] + n[138]);
p[47] = div_2*(n[139] + n[140] - n[141]);
p[48] = div_2*(n[142] + n[143] + n[144]);
p[49] = div_2*(n[145] + n[146] - n[147]);
p[50] = div_2*(n[148] - n[149])         ;
p[51] = div_2*(n[150] - n[151])         ;
p[52] = div_2*(n[152] + n[153] + n[154]);
p[53] = div_2*(n[155] + n[156] - n[157]);
p[54] = div_2*(n[158] + n[159] + n[160]);
p[55] = div_2*(n[161] + n[162] - n[163]);
p[56] = div_2*(n[164] + n[165] + n[166]);
p[57] = div_2*(n[167] + n[168] - n[169]);
p[58] = div_2*(n[170] + n[171] + n[172]);
p[59] = div_2*(n[173] + n[174] - n[175]);
p[60] = div_2*(n[176] + n[177] + n[178]);
p[61] = div_2*(n[179] + n[180] - n[181]);
p[62] = div_2*(n[182] + n[183] + n[184]);
p[63] = div_2*(n[185] + n[186] - n[187]);
p[64] = div_2*(n[188] + n[189] + n[190]);
p[65] = div_2*(n[191] + n[192] - n[193]);
p[66] = div_2*(n[194] + n[195] + n[196]);
p[67] = div_2*(n[197] + n[198] - n[199]);
p[68] = div_2*(n[200] + n[201] + n[202]);
p[69] = div_2*(n[203] + n[204] - n[205]);
p[70] = div_2*(n[206] + n[207] + n[208]);
p[71] = div_2*(n[209] + n[210] - n[211]);
p[72] = div_2*(n[212] + n[213] + n[214]);
p[73] = div_2*(n[215] + n[216] - n[217]);
p[74] = div_2*(n[218] + n[219] + n[220]);
p[75] = div_2*(n[221] + n[222] - n[223]);
p[76] = div_2*(n[224] + n[225] + n[226]);
p[77] = div_2*(n[227] + n[228] - n[229]);
p[78] = div_2*(n[230] + n[231] + n[232]);
p[79] = div_2*(n[233] + n[234] - n[235]);
p[80] = div_2*(n[236] + n[237] + n[238]);
p[81] = div_2*(n[239] + n[240] - n[241]);
p[82] = div_2*(n[242] + n[243] + n[244]);
p[83] = div_2*(n[245] + n[246] - n[247]);
p[84] = div_2*(n[248] + n[249] + n[250]);
p[85] = div_2*(n[251] + n[252] - n[253]);
p[86] = div_2*(n[254] + n[255] + n[256]);
p[87] = div_2*(n[257] + n[258] - n[259]);
p[88] = div_2*(n[260] + n[261] + n[262]);
p[89] = div_2*(n[263] + n[264] - n[265]);
p[90] = div_2*(n[266] + n[267] + n[268]);
p[91] = div_2*(n[269] + n[270] - n[271]);
p[92] = div_2*(n[272] + n[273] + n[274]);
p[93] = div_2*(n[275] + n[276] - n[277]);
p[94] = div_2*(n[278] + n[279] + n[280]);
p[95] = div_2*(n[281] + n[282] - n[283]);
p[96] = div_2*(n[284] + n[285] + n[286]);
p[97] = div_2*(n[287] + n[288] - n[289]);
p[98] = div_2*(n[290] + n[291] + n[292]);
p[99] = div_2*(n[293] + n[294] - n[295]);


re_X_0 = p[0][15:0] ;
im_X_0 = p[1][15:0] ;
re_X_1 = p[2][15:0] ;
 im_X_1 = p[3][15:0];
re_X_2 = p[4][15:0] ;
 im_X_2 = p[5][15:0];
re_X_3 = p[6][15:0] ;
 im_X_3 = p[7][15:0];
re_X_4 = p[8][15:0] ;
 im_X_4 = p[9][15:0];
re_X_5 = p[10][15:0] ;
 im_X_5 = p[11][15:0];
re_X_6 = p[12][15:0] ;
 im_X_6 = p[13][15:0];
re_X_7 = p[14][15:0] ;
 im_X_7 = p[15][15:0];
re_X_8 = p[16][15:0] ;
 im_X_8 = p[17][15:0];
re_X_9 = p[18][15:0] ;
 im_X_9 = p[19][15:0];
re_X_10 = p[20][15:0] ;
 im_X_10 = p[21][15:0];
re_X_11 = p[22][15:0] ;
 im_X_11 = p[23][15:0];
re_X_12 = p[24][15:0] ;
 im_X_12 = p[25][15:0];
re_X_13 = p[26][15:0] ;
 im_X_13 = p[27][15:0];
re_X_14 = p[28][15:0] ;
 im_X_14 = p[29][15:0];
re_X_15 = p[30][15:0] ;
 im_X_15 = p[31][15:0];
re_X_16 = p[32][15:0] ;
 im_X_16 = p[33][15:0];
re_X_17 = p[34][15:0] ;
 im_X_17 = p[35][15:0];
re_X_18 = p[36][15:0] ;
 im_X_18 = p[37][15:0];
re_X_19 = p[38][15:0] ;
 im_X_19 = p[39][15:0];
re_X_20 = p[40][15:0] ;
 im_X_20 = p[41][15:0];
re_X_21 = p[42][15:0] ;
 im_X_21 = p[43][15:0];
re_X_22 = p[44][15:0] ;
 im_X_22 = p[45][15:0];
re_X_23 = p[46][15:0] ;
 im_X_23 = p[47][15:0];
re_X_24 = p[48][15:0] ;
 im_X_24 = p[49][15:0];
re_X_25 = p[50][15:0] ;
 im_X_25 = p[51][15:0];
re_X_26 = p[52][15:0] ;
 im_X_26 = p[53][15:0];
re_X_27 = p[54][15:0] ;
 im_X_27 = p[55][15:0];
re_X_28 = p[56][15:0] ;
 im_X_28 = p[57][15:0];
re_X_29 = p[58][15:0] ;
 im_X_29 = p[59][15:0];
re_X_30 = p[60][15:0] ;
 im_X_30 = p[61][15:0];
re_X_31 = p[62][15:0] ;
 im_X_31 = p[63][15:0];
re_X_32 = p[64][15:0] ;
 im_X_32 = p[65][15:0];
re_X_33 = p[66][15:0] ;
 im_X_33 = p[67][15:0];
re_X_34 = p[68][15:0] ;
 im_X_34 = p[69][15:0];
re_X_35 = p[70][15:0] ;
 im_X_35 = p[71][15:0];
re_X_36 = p[72][15:0] ;
 im_X_36 = p[73][15:0];
re_X_37 = p[74][15:0] ;
 im_X_37 = p[75][15:0];
re_X_38 = p[76][15:0] ;
 im_X_38 = p[77][15:0];
re_X_39 = p[78][15:0] ;
 im_X_39 = p[79][15:0];
re_X_40 = p[80][15:0] ;
 im_X_40 = p[81][15:0];
re_X_41 = p[82][15:0] ;
 im_X_41 = p[83][15:0];
re_X_42 = p[84][15:0] ;
 im_X_42 = p[85][15:0];
re_X_43 = p[86][15:0] ;
 im_X_43 = p[87][15:0];
re_X_44 = p[88][15:0] ;
 im_X_44 = p[89][15:0];
re_X_45 = p[90][15:0] ;
 im_X_45 = p[91][15:0];
re_X_46 = p[92][15:0] ;
 im_X_46 = p[93][15:0];
re_X_47 = p[94][15:0] ;
 im_X_47 = p[95][15:0];
re_X_48 = p[96][15:0] ;
 im_X_48 = p[97][15:0];
re_X_49 = p[98][15:0] ;
 im_X_49 = p[99][15:0];

end

endmodule


///////////////////RADIX-5 1ST//////////////////////////////////////////////

module fft_radix5(clk,x11_r_0,x11_r_1,x11_r_2,x11_r_3,x11_r_4,x11_i_0,x11_i_1,x11_i_2,x11_i_3,x11_i_4,re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4);
input signed [15:0]x11_r_0,x11_r_1,x11_r_2,x11_r_3,x11_r_4,x11_i_0,x11_i_1,x11_i_2,x11_i_3,x11_i_4;
output reg signed [16:0]re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4;
wire signed [14:0]p_cos_36,n_cos_36,p_cos_72,n_cos_72,p_cos_0,n_sin_36,p_sin_36,p_sin_72,n_sin_72,div_5;
real p_cos_36_fract,n_cos_72_fract;
reg signed [30:0] z [81:0];
reg signed [15:0] y [81:0];
reg signed [31:0] m [9:0] ;
input clk;

assign p_cos_36='b011001111000110;
assign n_cos_36='b100110000111010;
assign p_cos_72='b001001111000110;
assign n_cos_72='b110110000111010;
assign p_cos_0= 'b011111111111111;
assign p_sin_36='b010010110011110;
assign n_sin_36='b101101001100010;
assign p_sin_72='b011110011011110;
assign n_sin_72='b100001100100010;
assign div_5   ='b000110011001100;
//////////////////////////////////////////// //output of re_X11_0

always@(posedge clk)
begin

z[9]= (x11_r_0 * p_cos_0 );
z[10]= (x11_r_1 * p_cos_0 );
z[11]= (x11_r_2 * p_cos_0 );
z[12]= (x11_r_3 * p_cos_0 );
z[13]= (x11_r_4 * p_cos_0 );

y[9] = z[9][30:15] + z[9][14];
y[10] = z[10][30:15] + z[10][14];
y[11] = z[11][30:15] + z[11][14];
y[12] = z[12][30:15] + z[12][14];
y[13] = z[13][30:15] + z[13][14];

///////////////////////////////////////////// //output of im_X11_0

z[14]= (x11_i_0 * p_cos_0 );
z[15]= (x11_i_1 * p_cos_0 );
z[16]= (x11_i_2 * p_cos_0 );
z[17]= (x11_i_3 * p_cos_0 );
z[18]= (x11_i_4 * p_cos_0 );

y[14] = z[14][30:15] + z[14][14];
y[15] = z[15][30:15] + z[15][14];
y[16] = z[16][30:15] + z[16][14];
y[17] = z[17][30:15] + z[17][14];
y[18] = z[18][30:15] + z[18][14];

////////////////////////////////////////////    //output of re_X11_1

z[0]= (x11_r_0 * p_cos_0);
z[1]= (x11_r_1 * p_cos_72);
z[2]= (x11_r_2 * n_cos_36);
z[3]= (x11_r_3 * n_cos_36);         
z[4]= (x11_r_4 * p_cos_72);
z[5]= (x11_i_1 * p_sin_72);
z[6]= (x11_i_2 * p_sin_36);
z[7]= (x11_i_3 * n_sin_36);
z[8]= (x11_i_4 * n_sin_72);

y[0] = z[0][30:15] + z[0][14];
y[1] = z[1][30:15] + z[1][14];
y[2] = z[2][30:15] + z[2][14];
y[3] = z[3][30:15] + z[3][14];
y[4] = z[4][30:15] + z[4][14];
y[5] = z[5][30:15] + z[5][14];
y[6] = z[6][30:15] + z[6][14];
y[7] = z[7][30:15] + z[7][14];
y[8] = z[8][30:15] + z[8][14];

/////////////////////////////////////////// //output of im_X11_1

z[19]= (x11_r_1 * p_sin_72);
z[20]= (x11_r_2 * p_sin_36);
z[21]= (x11_r_3 * n_sin_36);         
z[22]= (x11_r_4 * n_sin_72);
z[23]= (x11_i_0 * p_cos_0) ;
z[24]= (x11_i_1 * p_cos_72);
z[25]= (x11_i_2 * n_cos_36);
z[26]= (x11_i_3 * n_cos_36);
z[27]= (x11_i_4 * p_cos_72);

y[19] = z[19][30:15] + z[19][14];
y[20] = z[20][30:15] + z[20][14];
y[21] = z[21][30:15] + z[21][14];
y[22] = z[22][30:15] + z[22][14];
y[23] = z[23][30:15] + z[23][14];
y[24] = z[24][30:15] + z[24][14];
y[25] = z[25][30:15] + z[25][14];
y[26] = z[26][30:15] + z[26][14];
y[27] = z[27][30:15] + z[27][14];



/////////////////////////////////////////////output of re_X11_2

z[28]= (x11_r_0 * p_cos_0);
z[29]= (x11_r_1 * n_cos_36);
z[30]= (x11_r_2 * p_cos_72);
z[31]= (x11_r_3 * p_cos_72);         
z[32]= (x11_r_4 * n_cos_36);
z[33]= (x11_i_1 * p_sin_36);
z[34]= (x11_i_2 * n_sin_72);
z[35]= (x11_i_3 * p_sin_72);
z[36]= (x11_i_4 * n_sin_36);

y[28] = z[28][30:15] + z[28][14];
y[29] = z[29][30:15] + z[29][14];
y[30] = z[30][30:15] + z[30][14];
y[31] = z[31][30:15] + z[31][14];
y[32] = z[32][30:15] + z[32][14];
y[33] = z[33][30:15] + z[33][14];
y[34] = z[34][30:15] + z[34][14];
y[35] = z[35][30:15] + z[35][14];
y[36] = z[36][30:15] + z[36][14];

//////////////////////////////////////////////output of im_X11_2

z[37]= (x11_r_1 * p_sin_36);
z[38]= (x11_r_2 * n_sin_72);
z[39]= (x11_r_3 * p_sin_72);         
z[40]= (x11_r_4 * n_sin_36);
z[41]= (x11_i_0 * p_cos_0) ;
z[42]= (x11_i_1 * n_cos_36);
z[43]= (x11_i_2 * p_cos_72);
z[44]= (x11_i_3 * p_cos_72);
z[45]= (x11_i_4 * n_cos_36);

y[37]= z[37][30:15] + z[37][14]; 
y[38]= z[38][30:15] + z[38][14]; 
y[39]= z[39][30:15] + z[39][14];
y[40]= z[40][30:15] + z[40][14]; 
y[41]= z[41][30:15] + z[41][14]; 
y[42]= z[42][30:15] + z[42][14]; 
y[43]= z[43][30:15] + z[43][14]; 
y[44]= z[44][30:15] + z[44][14]; 
y[45]= z[45][30:15] + z[45][14];

////////////////////////////////////////////output of re_X11_3

z[46]= (x11_r_0 * p_cos_0);
z[47]= (x11_r_1 * n_cos_36);
z[48]= (x11_r_2 * p_cos_72);
z[49]= (x11_r_3 * p_cos_72);         
z[50]= (x11_r_4 * n_cos_36);
z[51]= (x11_i_1 * n_sin_36);
z[52]= (x11_i_2 * p_sin_72);
z[53]= (x11_i_3 * n_sin_72);
z[54]= (x11_i_4 * p_sin_36);

y[46]= z[46][30:15] + z[46][14]; 
y[47]= z[47][30:15] + z[47][14]; 
y[48]= z[48][30:15] + z[48][14]; 
y[49]= z[49][30:15] + z[49][14]; 
y[50]= z[50][30:15] + z[50][14]; 
y[51]= z[51][30:15] + z[51][14]; 
y[52]= z[52][30:15] + z[52][14]; 
y[53]= z[53][30:15] + z[53][14]; 
y[54]= z[54][30:15] + z[54][14];


///////////////////////////////////////////output of im_X11_3

z[55]= (x11_r_1 * n_sin_36);
z[56]= (x11_r_2 * p_sin_72);
z[57]= (x11_r_3 * n_sin_72);         
z[58]= (x11_r_4 * p_sin_36);
z[59]= (x11_i_0 * p_cos_0) ;
z[60]= (x11_i_1 * n_cos_36);
z[61]= (x11_i_2 * p_cos_72);
z[62]= (x11_i_3 * p_cos_72);
z[63]= (x11_i_4 * n_cos_36);

y[55]= z[55][30:15] + z[55][14]; 
y[56]= z[56][30:15] + z[56][14]; 
y[57]= z[57][30:15] + z[57][14]; 
y[58]= z[58][30:15] + z[58][14]; 
y[59]= z[59][30:15] + z[59][14]; 
y[60]= z[60][30:15] + z[60][14]; 
y[61]= z[61][30:15] + z[61][14]; 
y[62]= z[62][30:15] + z[62][14]; 
y[63]= z[63][30:15] + z[63][14];

////////////////////////////////////////////output of re_X11_4

z[64]= (x11_r_0 * p_cos_0);
z[65]= (x11_r_1 * p_cos_72);
z[66]= (x11_r_2 * n_cos_36);
z[67]= (x11_r_3 * n_cos_36);         
z[68]= (x11_r_4 * p_cos_72);
z[69]= (x11_i_1 * n_sin_72);
z[70]= (x11_i_2 * n_sin_36);
z[71]= (x11_i_3 * p_sin_36);
z[72]= (x11_i_4 * p_sin_72);

y[64]= z[64][30:15] + z[64][14]; 
y[65]= z[65][30:15] + z[65][14]; 
y[66]= z[66][30:15] + z[66][14]; 
y[67]= z[67][30:15] + z[67][14]; 
y[68]= z[68][30:15] + z[68][14]; 
y[69]= z[69][30:15] + z[69][14]; 
y[70]= z[70][30:15] + z[70][14]; 
y[71]= z[71][30:15] + z[71][14]; 
y[72]= z[72][30:15] + z[72][14];


///////////////////////////////////////////output of im_X11_4

z[73]= (x11_r_1 * n_sin_72);
z[74]= (x11_r_2 * n_sin_36);
z[75]= (x11_r_3 * p_sin_36);         
z[76]= (x11_r_4 * p_sin_72);
z[77]= (x11_i_0 * p_cos_0) ;
z[78]= (x11_i_1 * p_cos_72);
z[79]= (x11_i_2 * n_cos_36);
z[80]= (x11_i_3 * n_cos_36);
z[81]= (x11_i_4 * p_cos_72);

y[73]= z[73][30:15] + z[73][14]; 
y[74]= z[74][30:15] + z[74][14]; 
y[75]= z[75][30:15] + z[75][14]; 
y[76]= z[76][30:15] + z[76][14]; 
y[77]= z[77][30:15] + z[77][14]; 
y[78]= z[78][30:15] + z[78][14]; 
y[79]= z[79][30:15] + z[79][14]; 
y[80]= z[80][30:15] + z[80][14]; 
y[81]= z[81][30:15] + z[81][14];


/////////////////////////////////////////////


m[0] = div_5*(y[14] + y[15] + y[16] + y[17] + y[18]);
m[1] = div_5*(y[9]  + y[10] + y[11] + y[12] + y[13]);
m[2] = div_5*(y[0] + y[1] + y[2] + y[3] + y[4] + y[5] + y[6] + y[7] + y[8]);
m[3] = div_5*(y[23] - y[19] + y[24] - y[20] + y[25] - y[21] + y[26] - y[22] + y[27]);
m[4] = div_5*(y[28] + y[29] + y[30] + y[31] + y[32] + y[33] + y[34] + y[35] + y[36]);
m[5] = div_5*(y[41] - y[37] + y[42] - y[38] + y[43] - y[39] + y[44] - y[40] + y[45]);
m[6] = div_5*(y[46] + y[47] + y[48] + y[49] + y[50] + y[51] + y[52] + y[53] + y[54]);
m[7] = div_5*(y[59] - y[55] + y[60] - y[56] + y[61] - y[57] + y[62] - y[58] + y[63]);
m[8] = div_5*(y[64] + y[65] + y[66] + y[67] + y[68] + y[69] + y[70] + y[71] + y[72]);
m[9] = div_5*(y[77] - y[73] + y[78] - y[74] + y[79] - y[75] + y[80] - y[76] + y[81]);

im_X11_0 = m[0][28:12] + m[0][11] ;
re_X11_0 = m[1][28:12] + m[1][11] ;
im_X11_1 = m[3][28:12] + m[3][11] ;
re_X11_1 = m[2][28:12] + m[2][11] ;
im_X11_2 = m[5][28:12] + m[5][11] ;
re_X11_2 = m[4][28:12] + m[4][11] ;
im_X11_3 = m[7][28:12] + m[7][11] ;
re_X11_3 = m[6][28:12] + m[6][11] ;
im_X11_4 = m[9][28:12] + m[9][11] ;
re_X11_4 = m[8][28:12] + m[8][11] ;


end


endmodule


//////////////////RADIX-5 2ND//////////////////////////////////////////////////////////////////////////////////////


module radix_5_stage_2(clk,re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4,re_X12_0,im_X12_0,re_X12_1,im_X12_1,re_X12_2,im_X12_2,re_X12_3,im_X12_3,
re_X12_4,im_X12_4,re_X13_0,im_X13_0,re_X13_1,im_X13_1,re_X13_2,im_X13_2,re_X13_3,im_X13_3,re_X13_4,im_X13_4,re_X14_0,im_X14_0,re_X14_1,im_X14_1,re_X14_2,im_X14_2,re_X14_3,im_X14_3,
re_X14_4,im_X14_4,re_X15_0,im_X15_0,re_X15_1,im_X15_1,re_X15_2,im_X15_2,re_X15_3,im_X15_3,re_X15_4,im_X15_4,re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,
re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,
re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24);

input signed [16:0] re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4,re_X12_0,im_X12_0,re_X12_1,im_X12_1,re_X12_2,im_X12_2,re_X12_3,im_X12_3,
re_X12_4,im_X12_4,re_X13_0,im_X13_0,re_X13_1,im_X13_1,re_X13_2,im_X13_2,re_X13_3,im_X13_3,re_X13_4,im_X13_4,re_X14_0,im_X14_0,re_X14_1,im_X14_1,re_X14_2,im_X14_2,re_X14_3,im_X14_3,
re_X14_4,im_X14_4,re_X15_0,im_X15_0,re_X15_1,im_X15_1,re_X15_2,im_X15_2,re_X15_3,im_X15_3,re_X15_4,im_X15_4;

output reg signed [16:0] re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,
im_X1_8,re_X1_9,im_X1_9,re_X1_10,im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,re_X1_16,im_X1_16,re_X1_17,
im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24;

reg signed [31:0] q [441:0] ;
reg signed [15:0] p [441:0] ;
reg signed [31:0] m [49:0]  ;

input clk;

wire signed [14:0] p_cos_0,p_cos_14_4,p_sin_14_4,p_cos_28_8,p_sin_28_8,p_cos_43_2,p_sin_43_2,p_cos_57_6,p_sin_57_6,p_cos_72,p_sin_72,p_cos_86_4,p_sin_86_4,p_cos_100_8,p_sin_100_8,p_cos_115_2,
p_sin_115_2,p_cos_129_6,p_sin_129_6,p_cos_144,p_sin_144,p_cos_158_4,p_sin_158_4,p_cos_172_8,p_sin_172_8,p_cos_187_2,p_sin_187_2,p_cos_201_6,p_sin_201_6,p_cos_216,p_sin_216,p_cos_230_4,p_sin_230_4,
p_cos_244_8,p_sin_244_8,p_cos_259_2,p_sin_259_2,p_cos_273_6,p_sin_273_6,p_cos_288,p_sin_288,p_cos_302_4,p_sin_302_4,p_cos_316_8,p_sin_316_8,p_cos_331_2,p_sin_331_2,p_cos_345_6,p_sin_345_6,div_5;









assign p_cos_0     = 'b011111111111111;
assign p_cos_14_4  = 'b011110111111101;
assign p_sin_14_4  = 'b000111111101010;
assign p_cos_28_8  = 'b011100000010101;
assign p_sin_28_8  = 'b001111011010101;
assign p_cos_43_2  = 'b010111010100111;
assign p_sin_43_2  = 'b010101111001111;
assign p_cos_57_6  = 'b010001001001010;
assign p_sin_57_6  = 'b011011000001001;
assign p_cos_72    = 'b001001111000110;
assign p_sin_72    = 'b011110011011110;
assign p_cos_86_4  = 'b000010000000100;
assign p_sin_86_4  = 'b011111111011111;
assign p_cos_100_8 = 'b111010000000100;
assign p_sin_100_8 = 'b011111011011100;
assign p_cos_115_2 = 'b110010011000010;
assign p_sin_115_2 = 'b011100111101000;
assign p_cos_129_6 = 'b101011100110101;
assign p_sin_129_6 = 'b011000101001111;
assign p_cos_144   = 'b100110000111010;
assign p_sin_144   = 'b010010110011110;
assign p_cos_158_4 = 'b100010010000000;
assign p_sin_158_4 = 'b001011110001110;
assign p_cos_172_8 = 'b100000010000010;
assign p_sin_172_8 = 'b000100000000101;
assign p_cos_187_2 = 'b100000010000010;
assign p_sin_187_2 = 'b111011111111011;
assign p_cos_201_6 = 'b100010010000000;
assign p_sin_201_6 = 'b110100001110010;
assign p_cos_216   = 'b100110000111010;
assign p_sin_216   = 'b101101001100010;
assign p_cos_230_4 = 'b101011100110101;
assign p_sin_230_4 = 'b100111010110001;
assign p_cos_244_8 = 'b110010011000010;
assign p_sin_244_8 = 'b100011000011000;
assign p_cos_259_2 = 'b111010000000100;
assign p_sin_259_2 = 'b100000100100100;
assign p_cos_273_6 = 'b000010000000100;
assign p_sin_273_6 = 'b100000000100001;
assign p_cos_288   = 'b001001111000110;
assign p_sin_288   = 'b100001100100010;
assign p_cos_302_4 = 'b010001001001010;
assign p_sin_302_4 = 'b100100111110111;
assign p_cos_316_8 = 'b010111010100111;
assign p_sin_316_8 = 'b101010000110001;
assign p_cos_331_2 = 'b011100000010101;
assign p_sin_331_2 = 'b110000100101011;
assign p_cos_345_6 = 'b011110111111101;
assign p_sin_345_6 = 'b111000000010110;
assign div_5   ='b000110011001100;


///////////////////////////////////////////////////////////////// output of re_X1_0

always@(posedge clk)
begin

q[0]= (re_X11_0 * p_cos_0 );
q[1]= (re_X12_0 * p_cos_0 );
q[2]= (re_X13_0 * p_cos_0 );
q[3]= (re_X14_0 * p_cos_0 );
q[4]= (re_X15_0 * p_cos_0 );

p[0] = q[0][31:16] + q[0][15];
p[1] = q[1][31:16] + q[1][15];
p[2] = q[2][31:16] + q[2][15];
p[3] = q[3][31:16] + q[3][15];
p[4] = q[4][31:16] + q[4][15];

////////////////////////////////////////////////////////////////////// output of im_X1_0

q[5]= (im_X11_0 * p_cos_0 );
q[6]= (im_X12_0 * p_cos_0 );
q[7]= (im_X13_0 * p_cos_0 );
q[8]= (im_X14_0 * p_cos_0 );
q[9]= (im_X15_0 * p_cos_0 );


p[5] = q[5][31:16] + q[5][15];
p[6] = q[6][31:16] + q[6][15];
p[7] = q[7][31:16] + q[7][15];
p[8] = q[8][31:16] + q[8][15];
p[9] = q[9][31:16] + q[9][15];

/////////////////////////////////////////////////////////////////////////////////// output of re_X1_1

q[10]= (re_X11_1 * p_cos_0 );
q[11]= (re_X12_1 * p_cos_14_4 );
q[12]= (re_X13_1 * p_cos_28_8 );
q[13]= (re_X14_1 * p_cos_43_2 );
q[14]= (re_X15_1 * p_cos_57_6 );
q[15]= (im_X12_1 * p_sin_14_4 );
q[16]= (im_X13_1 * p_sin_28_8 );
q[17]= (im_X14_1 * p_sin_43_2 );
q[18]= (im_X15_1 * p_sin_57_6 );

p[10] = q[10][31:16] + q[10][15];
p[11] = q[11][31:16] + q[11][15];
p[12] = q[12][31:16] + q[12][15];
p[13] = q[13][31:16] + q[13][15];
p[14] = q[14][31:16] + q[14][15];
p[15] = q[15][31:16] + q[15][15];
p[16] = q[16][31:16] + q[16][15];
p[17] = q[17][31:16] + q[17][15];
p[18] = q[18][31:16] + q[18][15];


////////////////////////////////////////////////////////////////////////////////// output of im_X1_1

q[19]= (im_X11_1 * p_cos_0 );
q[20]= (im_X12_1 * p_cos_14_4 );
q[21]= (im_X13_1 * p_cos_28_8 );
q[22]= (im_X14_1 * p_cos_43_2 );
q[23]= (im_X15_1 * p_cos_57_6 );
q[24]= (re_X12_1 * p_sin_14_4 );
q[25]= (re_X13_1 * p_sin_28_8 );
q[26]= (re_X14_1 * p_sin_43_2 );
q[27]= (re_X15_1 * p_sin_57_6 );

p[19] = q[19][31:16] + q[19][15];
p[20] = q[20][31:16] + q[20][15];
p[21] = q[21][31:16] + q[21][15];
p[22] = q[22][31:16] + q[22][15];
p[23] = q[23][31:16] + q[23][15];
p[24] = q[24][31:16] + q[24][15];
p[25] = q[25][31:16] + q[25][15];
p[26] = q[26][31:16] + q[26][15];
p[27] = q[27][31:16] + q[27][15];

/////////////////////////////////////////////////////////////////////////////////// output of re_X1_2

q[28]= (re_X11_2 * p_cos_0 );
q[29]= (re_X12_2 * p_cos_28_8 );
q[30]= (re_X13_2 * p_cos_57_6 );
q[31]= (re_X14_2 * p_cos_86_4 );
q[32]= (re_X15_2 * p_cos_115_2 );
q[33]= (im_X12_2 * p_sin_28_8 );
q[34]= (im_X13_2 * p_sin_57_6 );
q[35]= (im_X14_2 * p_sin_86_4 );
q[36]= (im_X15_2 * p_sin_115_2 );

p[28] = q[28][31:16] + q[28][15];
p[29] = q[29][31:16] + q[29][15];
p[30] = q[30][31:16] + q[30][15];
p[31] = q[31][31:16] + q[31][15];
p[32] = q[32][31:16] + q[32][15];
p[33] = q[33][31:16] + q[33][15];
p[34] = q[34][31:16] + q[34][15];
p[35] = q[35][31:16] + q[35][15];
p[36] = q[36][31:16] + q[36][15];

////////////////////////////////////////////////////////////////////////////////////// output of im_X1_2

q[37]= (im_X11_2 * p_cos_0 );
q[38]= (im_X12_2 * p_cos_28_8 );
q[39]= (im_X13_2 * p_cos_57_6 );
q[40]= (im_X14_2 * p_cos_86_4 );
q[41]= (im_X15_2 * p_cos_115_2 );
q[42]= (re_X12_2 * p_sin_28_8 );
q[43]= (re_X13_2 * p_sin_57_6 );
q[44]= (re_X14_2 * p_sin_86_4 );
q[45]= (re_X15_2 * p_sin_115_2 );

p[37] = q[37][31:16] + q[37][15];
p[38] = q[38][31:16] + q[38][15];
p[39] = q[39][31:16] + q[39][15];
p[40] = q[40][31:16] + q[40][15];
p[41] = q[41][31:16] + q[41][15];
p[42] = q[42][31:16] + q[42][15];
p[43] = q[43][31:16] + q[43][15];
p[44] = q[44][31:16] + q[44][15];
p[45] = q[45][31:16] + q[45][15];

/////////////////////////////////////////////////////////////////////////////////////// output of re_X1_3

q[46]= (re_X11_3 * p_cos_0 );
q[47]= (re_X12_3 * p_cos_43_2 );
q[48]= (re_X13_3 * p_cos_86_4 );
q[49]= (re_X14_3 * p_cos_129_6 );
q[50]= (re_X15_3 * p_cos_172_8 );
q[51]= (im_X12_3 * p_sin_43_2 );
q[52]= (im_X13_3 * p_sin_86_4 );
q[53]= (im_X14_3 * p_sin_129_6 );
q[54]= (im_X15_3 * p_sin_172_8 );

p[46] = q[46][31:16] + q[46][15];
p[47] = q[47][31:16] + q[47][15];
p[48] = q[48][31:16] + q[48][15];
p[49] = q[49][31:16] + q[49][15];
p[50] = q[50][31:16] + q[50][15];
p[51] = q[51][31:16] + q[51][15];
p[52] = q[52][31:16] + q[52][15];
p[53] = q[53][31:16] + q[53][15];
p[54] = q[54][31:16] + q[54][15];

////////////////////////////////////////////////////////////////////////////////////// output of im_X1_3

q[55]= (im_X11_3 * p_cos_0 );
q[56]= (im_X12_3 * p_cos_43_2 );
q[57]= (im_X13_3 * p_cos_86_4 );
q[58]= (im_X14_3 * p_cos_129_6 );
q[59]= (im_X15_3 * p_cos_172_8 );
q[60]= (re_X12_3 * p_sin_43_2 );
q[61]= (re_X13_3 * p_sin_86_4 );
q[62]= (re_X14_3 * p_sin_129_6 );
q[63]= (re_X15_3 * p_sin_172_8 );

p[55] = q[55][31:16] + q[55][15];
p[56] = q[56][31:16] + q[56][15];
p[57] = q[57][31:16] + q[57][15];
p[58] = q[58][31:16] + q[58][15];
p[59] = q[59][31:16] + q[59][15];
p[60] = q[60][31:16] + q[60][15];
p[61] = q[61][31:16] + q[61][15];
p[62] = q[62][31:16] + q[62][15];
p[63] = q[63][31:16] + q[63][15];

////////////////////////////////////////////////////////////////////////////////////// output of re_X1_4

q[64]= (re_X11_4 * p_cos_0 );
q[65]= (re_X12_4 * p_cos_57_6 );
q[66]= (re_X13_4 * p_cos_115_2 );
q[67]= (re_X14_4 * p_cos_172_8 );
q[68]= (re_X15_4 * p_cos_230_4 );
q[69]= (im_X12_4 * p_sin_57_6 );
q[70]= (im_X13_4 * p_sin_115_2 );
q[71]= (im_X14_4 * p_sin_172_8 );
q[72]= (im_X15_4 * p_sin_230_4 );

p[64] = q[64][31:16] + q[64][15];
p[65] = q[65][31:16] + q[65][15];
p[66] = q[66][31:16] + q[66][15];
p[67] = q[67][31:16] + q[67][15];
p[68] = q[68][31:16] + q[68][15];
p[69] = q[69][31:16] + q[69][15];
p[70] = q[70][31:16] + q[70][15];
p[71] = q[71][31:16] + q[71][15];
p[72] = q[72][31:16] + q[72][15];


//////////////////////////////////////////////////////////////////////////////////////// output of im_X1_4

q[73]= (im_X11_4 * p_cos_0 );
q[74]= (im_X12_4 * p_cos_57_6 );
q[75]= (im_X13_4 * p_cos_115_2 );
q[76]= (im_X14_4 * p_cos_172_8 );
q[77]= (im_X15_4 * p_cos_230_4 );
q[78]= (re_X12_4 * p_sin_57_6 );
q[79]= (re_X13_4 * p_sin_115_2 );
q[80]= (re_X14_4 * p_sin_172_8 );
q[81]= (re_X15_4 * p_sin_230_4 );
 
p[73] = q[73][31:16] + q[73][15];
p[74] = q[74][31:16] + q[74][15];
p[75] = q[75][31:16] + q[75][15];
p[76] = q[76][31:16] + q[76][15];
p[77] = q[77][31:16] + q[77][15];
p[78] = q[78][31:16] + q[78][15];
p[79] = q[79][31:16] + q[79][15];
p[80] = q[80][31:16] + q[80][15];
p[81] = q[81][31:16] + q[81][15];

////////////////////////////////////////////////////////////////////////////////////// output of re_X1_5

q[82]= (re_X11_0 * p_cos_0 );
q[83]= (re_X12_0 * p_cos_72 );
q[84]= (re_X13_0 * p_cos_144 );
q[85]= (re_X14_0 * p_cos_216 );
q[86]= (re_X15_0 * p_cos_288 );
q[87]= (im_X12_0 * p_sin_72 );
q[88]= (im_X13_0 * p_sin_144 );
q[89]= (im_X14_0 * p_sin_216 );
q[90]= (im_X15_0 * p_sin_288 );

p[82] = q[82][31:16] + q[82][15];
p[83] = q[83][31:16] + q[83][15];
p[84] = q[84][31:16] + q[84][15];
p[85] = q[85][31:16] + q[85][15];
p[86] = q[86][31:16] + q[86][15];
p[87] = q[87][31:16] + q[87][15];
p[88] = q[88][31:16] + q[88][15];
p[89] = q[89][31:16] + q[89][15];
p[90] = q[90][31:16] + q[90][15];

////////////////////////////////////////////////////////////////////////////////////// output of im_X1_5

q[91]= (im_X11_0 * p_cos_0 );
q[92]= (im_X12_0 * p_cos_72 );
q[93]= (im_X13_0 * p_cos_144 );
q[94]= (im_X14_0 * p_cos_216 );
q[95]= (im_X15_0 * p_cos_288 );
q[96]= (re_X12_0 * p_sin_72 );
q[97]= (re_X13_0 * p_sin_144 );
q[98]= (re_X14_0 * p_sin_216 );
q[99]= (re_X15_0 * p_sin_288 );

p[91] = q[91][31:16] + q[91][15];
p[92] = q[92][31:16] + q[92][15];
p[93] = q[93][31:16] + q[93][15];
p[94] = q[94][31:16] + q[94][15];
p[95] = q[95][31:16] + q[95][15];
p[96] = q[96][31:16] + q[96][15];
p[97] = q[97][31:16] + q[97][15];
p[98] = q[98][31:16] + q[98][15];
p[99] = q[99][31:16] + q[99][15];

//////////////////////////////////////////////////////////////////////////////////////// output of re_X1_6

q[100]= (re_X11_1 * p_cos_0 );
q[101]= (re_X12_1 * p_cos_86_4 );
q[102]= (re_X13_1 * p_cos_172_8 );
q[103]= (re_X14_1 * p_cos_259_2 );
q[104]= (re_X15_1 * p_cos_345_6 );
q[105]= (im_X12_1 * p_sin_86_4 );
q[106]= (im_X13_1 * p_sin_172_8 );
q[107]= (im_X14_1 * p_sin_259_2 );
q[108]= (im_X15_1 * p_sin_345_6 );

p[100] = q[100][31:16] + q[100][15];
p[101] = q[101][31:16] + q[101][15];
p[102] = q[102][31:16] + q[102][15];
p[103] = q[103][31:16] + q[103][15];
p[104] = q[104][31:16] + q[104][15];
p[105] = q[105][31:16] + q[105][15];
p[106] = q[106][31:16] + q[106][15];
p[107] = q[107][31:16] + q[107][15];
p[108] = q[108][31:16] + q[108][15];

//////////////////////////////////////////////////////////////////////////////////////// output of im_X1_6

q[109]= (im_X11_1 * p_cos_0 );
q[110]= (im_X12_1 * p_cos_86_4 );
q[111]= (im_X13_1 * p_cos_172_8 );
q[112]= (im_X14_1 * p_cos_259_2 );
q[113]= (im_X15_1 * p_cos_345_6 );
q[114]= (re_X12_1 * p_sin_86_4 );
q[115]= (re_X13_1 * p_sin_172_8 );
q[116]= (re_X14_1 * p_sin_259_2 );
q[117]= (re_X15_1 * p_sin_345_6 );

p[109] = q[109][31:16] + q[109][15];
p[110] = q[110][31:16] + q[110][15];
p[111] = q[111][31:16] + q[111][15];
p[112] = q[112][31:16] + q[112][15];
p[113] = q[113][31:16] + q[113][15];
p[114] = q[114][31:16] + q[114][15];
p[115] = q[115][31:16] + q[115][15];
p[116] = q[116][31:16] + q[116][15];
p[117] = q[117][31:16] + q[117][15];

//////////////////////////////////////////////////////////////////////////////////////// output of re_X1_7

q[118]= (re_X11_2 * p_cos_0 );
q[119]= (re_X12_2 * p_cos_100_8 );
q[120]= (re_X13_2 * p_cos_201_6 );
q[121]= (re_X14_2 * p_cos_302_4 );
q[122]= (re_X15_2 * p_cos_43_2 );
q[123]= (im_X12_2 * p_sin_100_8 );
q[124]= (im_X13_2 * p_sin_201_6 );
q[125]= (im_X14_2 * p_sin_302_4 );
q[126]= (im_X15_2 * p_sin_43_2 );

p[118] = q[118][31:16] + q[118][15];
p[119] = q[119][31:16] + q[119][15];
p[120] = q[120][31:16] + q[120][15];
p[121] = q[121][31:16] + q[121][15];
p[122] = q[122][31:16] + q[122][15];
p[123] = q[123][31:16] + q[123][15];
p[124] = q[124][31:16] + q[124][15];
p[125] = q[125][31:16] + q[125][15];
p[126] = q[126][31:16] + q[126][15];

/////////////////////////////////////////////////////////////////////////////////////// output of im_X1_7

q[127]= (im_X11_2 * p_cos_0 );
q[128]= (im_X12_2 * p_cos_100_8 );
q[129]= (im_X13_2 * p_cos_201_6 );
q[130]= (im_X14_2 * p_cos_302_4 );
q[131]= (im_X15_2 * p_cos_43_2 );
q[132]= (re_X12_2 * p_sin_100_8 );
q[133]= (re_X13_2 * p_sin_201_6 );
q[134]= (re_X14_2 * p_sin_302_4 );
q[135]= (re_X15_2 * p_sin_43_2 );

p[127] = q[127][31:16] + q[127][15];
p[128] = q[128][31:16] + q[128][15];
p[129] = q[129][31:16] + q[129][15];
p[130] = q[130][31:16] + q[130][15];
p[131] = q[131][31:16] + q[131][15];
p[132] = q[132][31:16] + q[132][15];
p[133] = q[133][31:16] + q[133][15];
p[134] = q[134][31:16] + q[134][15];
p[135] = q[135][31:16] + q[135][15];

///////////////////////////////////////////////////////////////////////////////////// output of re_X1_8

q[136]= (re_X11_3 * p_cos_0 );
q[137]= (re_X12_3 * p_cos_115_2 );
q[138]= (re_X13_3 * p_cos_230_4 );
q[139]= (re_X14_3 * p_cos_345_6 );
q[140]= (re_X15_3 * p_cos_100_8 );
q[141]= (im_X12_3 * p_sin_115_2 );
q[142]= (im_X13_3 * p_sin_230_4 );
q[143]= (im_X14_3 * p_sin_345_6 );
q[144]= (im_X15_3 * p_sin_100_8 );

p[136] = q[136][31:16] + q[136][15];
p[137] = q[137][31:16] + q[137][15];
p[138] = q[138][31:16] + q[138][15];
p[139] = q[139][31:16] + q[139][15];
p[140] = q[140][31:16] + q[140][15];
p[141] = q[141][31:16] + q[141][15];
p[142] = q[142][31:16] + q[142][15];
p[143] = q[143][31:16] + q[143][15];
p[144] = q[144][31:16] + q[144][15];

///////////////////////////////////////////////////////////////////////////////////// output of im_X1_8

q[145]= (im_X11_3 * p_cos_0 );
q[146]= (im_X12_3 * p_cos_115_2 );
q[147]= (im_X13_3 * p_cos_230_4 );
q[148]= (im_X14_3 * p_cos_345_6 );
q[149]= (im_X15_3 * p_cos_100_8 );
q[150]= (re_X12_3 * p_sin_115_2 );
q[151]= (re_X13_3 * p_sin_230_4 );
q[152]= (re_X14_3 * p_sin_345_6 );
q[153]= (re_X15_3 * p_sin_100_8 );

p[145] = q[145][31:16] + q[145][15];
p[146] = q[146][31:16] + q[146][15];
p[147] = q[147][31:16] + q[147][15];
p[148] = q[148][31:16] + q[148][15];
p[149] = q[149][31:16] + q[149][15];
p[150] = q[150][31:16] + q[150][15];
p[151] = q[151][31:16] + q[151][15];
p[152] = q[152][31:16] + q[152][15];
p[153] = q[153][31:16] + q[153][15];

/////////////////////////////////////////////////////////////////////////////////////// output of re_X1_9

q[154]= (re_X11_4 * p_cos_0 );
q[155]= (re_X12_4 * p_cos_129_6 );
q[156]= (re_X13_4 * p_cos_259_2 );
q[157]= (re_X14_4 * p_cos_28_8 );
q[158]= (re_X15_4 * p_cos_158_4 );
q[159]= (im_X12_4 * p_sin_129_6 );
q[160]= (im_X13_4 * p_sin_259_2 );
q[161]= (im_X14_4 * p_sin_28_8 );
q[162]= (im_X15_4 * p_sin_158_4 );

p[154] = q[154][31:16] + q[154][15];
p[155] = q[155][31:16] + q[155][15];
p[156] = q[156][31:16] + q[156][15];
p[157] = q[157][31:16] + q[157][15];
p[158] = q[158][31:16] + q[158][15];
p[159] = q[159][31:16] + q[159][15];
p[160] = q[160][31:16] + q[160][15];
p[161] = q[161][31:16] + q[161][15];
p[162] = q[162][31:16] + q[162][15];


///////////////////////////////////////////////////////////////////////////////////// output of im_X1_9

q[163]= (im_X11_4 * p_cos_0 );
q[164]= (im_X12_4 * p_cos_129_6 );
q[165]= (im_X13_4 * p_cos_259_2 );
q[166]= (im_X14_4 * p_cos_28_8 );
q[167]= (im_X15_4 * p_cos_158_4 );
q[168]= (re_X12_4 * p_sin_129_6 );
q[169]= (re_X13_4 * p_sin_259_2 );
q[170]= (re_X14_4 * p_sin_28_8 );
q[171]= (re_X15_4 * p_sin_158_4 );

p[163] = q[163][31:16] + q[163][15];
p[164] = q[164][31:16] + q[164][15];
p[165] = q[165][31:16] + q[165][15];
p[166] = q[166][31:16] + q[166][15];
p[167] = q[167][31:16] + q[167][15];
p[168] = q[168][31:16] + q[168][15];
p[169] = q[169][31:16] + q[169][15];
p[170] = q[170][31:16] + q[170][15];
p[171] = q[171][31:16] + q[171][15];

///////////////////////////////////////////////////////////////////////////////////////// output of re_X1_10

q[172]= (re_X11_0 * p_cos_0 );
q[173]= (re_X12_0 * p_cos_144 );
q[174]= (re_X13_0 * p_cos_288 );
q[175]= (re_X14_0 * p_cos_72 );
q[176]= (re_X15_0 * p_cos_216 );
q[177]= (im_X12_0 * p_sin_144 );
q[178]= (im_X13_0 * p_sin_288 );
q[179]= (im_X14_0 * p_sin_72 );
q[180]= (im_X15_0 * p_sin_216 );

p[172] = q[172][31:16] + q[172][15];
p[173] = q[173][31:16] + q[173][15];
p[174] = q[174][31:16] + q[174][15];
p[175] = q[175][31:16] + q[175][15];
p[176] = q[176][31:16] + q[176][15];
p[177] = q[177][31:16] + q[177][15];
p[178] = q[178][31:16] + q[178][15];
p[179] = q[179][31:16] + q[179][15];
p[180] = q[180][31:16] + q[180][15];


////////////////////////////////////////////////////////////////////////////////////////// output of im_X1_10

q[181]= (im_X11_0 * p_cos_0 );
q[182]= (im_X12_0 * p_cos_144 );
q[183]= (im_X13_0 * p_cos_288 );
q[184]= (im_X14_0 * p_cos_72 );
q[185]= (im_X15_0 * p_cos_216 );
q[186]= (re_X12_0 * p_sin_144 );
q[187]= (re_X13_0 * p_sin_288 );
q[188]= (re_X14_0 * p_sin_72 );
q[189]= (re_X15_0 * p_sin_216 );

p[181] = q[181][31:16] + q[181][15];
p[182] = q[182][31:16] + q[182][15];
p[183] = q[183][31:16] + q[183][15];
p[184] = q[184][31:16] + q[184][15];
p[185] = q[185][31:16] + q[185][15];
p[186] = q[186][31:16] + q[186][15];
p[187] = q[187][31:16] + q[187][15];
p[188] = q[188][31:16] + q[188][15];
p[189] = q[189][31:16] + q[189][15];

/////////////////////////////////////////////////////////////////////////////////////// output of re_X1_11

q[190]= (re_X11_1 * p_cos_0 );
q[191]= (re_X12_1 * p_cos_158_4 );
q[192]= (re_X13_1 * p_cos_316_8 );
q[193]= (re_X14_1 * p_cos_115_2 );
q[194]= (re_X15_1 * p_cos_273_6 );
q[195]= (im_X12_1 * p_sin_158_4 );
q[196]= (im_X13_1 * p_sin_316_8 );
q[197]= (im_X14_1 * p_sin_115_2 );
q[198]= (im_X15_1 * p_sin_273_6 );

p[190] = q[190][31:16] + q[190][15];
p[191] = q[191][31:16] + q[191][15];
p[192] = q[192][31:16] + q[192][15];
p[193] = q[193][31:16] + q[193][15];
p[194] = q[194][31:16] + q[194][15];
p[195] = q[195][31:16] + q[195][15];
p[196] = q[196][31:16] + q[196][15];
p[197] = q[197][31:16] + q[197][15];
p[198] = q[198][31:16] + q[198][15];

//////////////////////////////////////////////////////////////////////////////////////// output of im_X1_11

q[199]= (im_X11_1 * p_cos_0 );
q[200]= (im_X12_1 * p_cos_158_4 );
q[201]= (im_X13_1 * p_cos_316_8 );
q[202]= (im_X14_1 * p_cos_115_2 );
q[203]= (im_X15_1 * p_cos_273_6 );
q[204]= (re_X12_1 * p_sin_158_4 );
q[205]= (re_X13_1 * p_sin_316_8 );
q[206]= (re_X14_1 * p_sin_115_2 );
q[207]= (re_X15_1 * p_sin_273_6 );

p[199] = q[199][31:16] + q[199][15];
p[200] = q[200][31:16] + q[200][15];
p[201] = q[201][31:16] + q[201][15];
p[202] = q[202][31:16] + q[202][15];
p[203] = q[203][31:16] + q[203][15];
p[204] = q[204][31:16] + q[204][15];
p[205] = q[205][31:16] + q[205][15];
p[206] = q[206][31:16] + q[206][15];
p[207] = q[207][31:16] + q[207][15];

///////////////////////////////////////////////////////////////////////////////////////// output of re_X1_12

q[208]= (re_X11_2 * p_cos_0 );
q[209]= (re_X12_2 * p_cos_172_8 );
q[210]= (re_X13_2 * p_cos_345_6 );
q[211]= (re_X14_2 * p_cos_158_4 );
q[212]= (re_X15_2 * p_cos_331_2 );
q[213]= (im_X12_2 * p_sin_172_8 );
q[214]= (im_X13_2 * p_sin_345_6 );
q[215]= (im_X14_2 * p_sin_158_4 );
q[216]= (im_X15_2 * p_sin_331_2 );

p[208] = q[208][31:16] + q[208][15];
p[209] = q[209][31:16] + q[209][15];
p[210] = q[210][31:16] + q[210][15];
p[211] = q[211][31:16] + q[211][15];
p[212] = q[212][31:16] + q[212][15];
p[213] = q[213][31:16] + q[213][15];
p[214] = q[214][31:16] + q[214][15];
p[215] = q[215][31:16] + q[215][15];
p[216] = q[216][31:16] + q[216][15];

//////////////////////////////////////////////////////////////////////////////////////// output of im_X1_12

q[217]= (im_X11_2 * p_cos_0 );
q[218]= (im_X12_2 * p_cos_172_8 );
q[219]= (im_X13_2 * p_cos_345_6 );
q[220]= (im_X14_2 * p_cos_158_4 );
q[221]= (im_X15_2 * p_cos_331_2 );
q[222]= (re_X12_2 * p_sin_172_8 );
q[223]= (re_X13_2 * p_sin_345_6 );
q[224]= (re_X14_2 * p_sin_158_4 );
q[225]= (re_X15_2 * p_sin_331_2 );

p[217] = q[217][31:16] + q[217][15];
p[218] = q[218][31:16] + q[218][15];
p[219] = q[219][31:16] + q[219][15];
p[220] = q[220][31:16] + q[220][15];
p[221] = q[221][31:16] + q[221][15];
p[222] = q[222][31:16] + q[222][15];
p[223] = q[223][31:16] + q[223][15];
p[224] = q[224][31:16] + q[224][15];
p[225] = q[225][31:16] + q[225][15];

/////////////////////////////////////////////////////////////////////////////////////// output of re_X1_13

q[226]= (re_X11_3 * p_cos_0 );
q[227]= (re_X12_3 * p_cos_187_2 );
q[228]= (re_X13_3 * p_cos_14_4 );
q[229]= (re_X14_3 * p_cos_201_6 );
q[230]= (re_X15_3 * p_cos_28_8 );
q[231]= (im_X12_3 * p_sin_187_2 );
q[232]= (im_X13_3 * p_sin_14_4 );
q[233]= (im_X14_3 * p_sin_201_6 );
q[234]= (im_X15_3 * p_sin_28_8 );

p[226] = q[226][31:16] + q[226][15];
p[227] = q[227][31:16] + q[227][15];
p[228] = q[228][31:16] + q[228][15];
p[229] = q[229][31:16] + q[229][15];
p[230] = q[230][31:16] + q[230][15];
p[231] = q[231][31:16] + q[231][15];
p[232] = q[232][31:16] + q[232][15];
p[233] = q[233][31:16] + q[233][15];
p[234] = q[234][31:16] + q[234][15];

/////////////////////////////////////////////////////////////////////////////////////// output of im_X1_13

q[235]= (im_X11_3 * p_cos_0 );
q[236]= (im_X12_3 * p_cos_187_2 );
q[237]= (im_X13_3 * p_cos_14_4 );
q[238]= (im_X14_3 * p_cos_201_6 );
q[239]= (im_X15_3 * p_cos_28_8 );
q[240]= (re_X12_3 * p_sin_187_2 );
q[241]= (re_X13_3 * p_sin_14_4 );
q[242]= (re_X14_3 * p_sin_201_6 );
q[243]= (re_X15_3 * p_sin_28_8 );

p[235] = q[235][31:16] + q[235][15];
p[236] = q[236][31:16] + q[236][15];
p[237] = q[237][31:16] + q[237][15];
p[238] = q[238][31:16] + q[238][15];
p[239] = q[239][31:16] + q[239][15];
p[240] = q[240][31:16] + q[240][15];
p[241] = q[241][31:16] + q[241][15];
p[242] = q[242][31:16] + q[242][15];
p[243] = q[243][31:16] + q[243][15];

//////////////////////////////////////////////////////////////////////////////////////// output of re_X1_14

q[244]= (re_X11_4 * p_cos_0 );
q[245]= (re_X12_4 * p_cos_201_6 );
q[246]= (re_X13_4 * p_cos_43_2 );
q[247]= (re_X14_4 * p_cos_244_8 );
q[248]= (re_X15_4 * p_cos_86_4 );
q[249]= (im_X12_4 * p_sin_201_6 );
q[250]= (im_X13_4 * p_sin_43_2 );
q[251]= (im_X14_4 * p_sin_244_8 );
q[252]= (im_X15_4 * p_sin_86_4 );

p[244] = q[244][31:16] + q[244][15];
p[245] = q[245][31:16] + q[245][15];
p[246] = q[246][31:16] + q[246][15];
p[247] = q[247][31:16] + q[247][15];
p[248] = q[248][31:16] + q[248][15];
p[249] = q[249][31:16] + q[249][15];
p[250] = q[250][31:16] + q[250][15];
p[251] = q[251][31:16] + q[251][15];
p[252] = q[252][31:16] + q[252][15];

///////////////////////////////////////////////////////////////////////////////////////// output of im_X1_14

q[253]= (im_X11_4 * p_cos_0 );
q[254]= (im_X12_4 * p_cos_201_6 );
q[255]= (im_X13_4 * p_cos_43_2 );
q[256]= (im_X14_4 * p_cos_244_8 );
q[257]= (im_X15_4 * p_cos_86_4 );
q[258]= (re_X12_4 * p_sin_201_6 );
q[259]= (re_X13_4 * p_sin_43_2 );
q[260]= (re_X14_4 * p_sin_244_8 );
q[261]= (re_X15_4 * p_sin_86_4 );

p[253] = q[253][31:16] + q[253][15];
p[254] = q[254][31:16] + q[254][15];
p[255] = q[255][31:16] + q[255][15];
p[256] = q[256][31:16] + q[256][15];
p[257] = q[257][31:16] + q[257][15];
p[258] = q[258][31:16] + q[258][15];
p[259] = q[259][31:16] + q[259][15];
p[260] = q[260][31:16] + q[260][15];
p[261] = q[261][31:16] + q[261][15];

///////////////////////////////////////////////////////////////////////////////////////// output of re_X1_15

q[262]= (re_X11_0 * p_cos_0 );
q[263]= (re_X12_0 * p_cos_216 );
q[264]= (re_X13_0 * p_cos_72 );
q[265]= (re_X14_0 * p_cos_288 );
q[266]= (re_X15_0 * p_cos_144 );
q[267]= (im_X12_0 * p_sin_216 );
q[268]= (im_X13_0 * p_sin_72 );
q[269]= (im_X14_0 * p_sin_288 );
q[270]= (im_X15_0 * p_sin_144 );

p[262] = q[262][31:16] + q[262][15];
p[263] = q[263][31:16] + q[263][15];
p[264] = q[264][31:16] + q[264][15];
p[265] = q[265][31:16] + q[265][15];
p[266] = q[266][31:16] + q[266][15];
p[267] = q[267][31:16] + q[267][15];
p[268] = q[268][31:16] + q[268][15];
p[269] = q[269][31:16] + q[269][15];

//////////////////////////////////////////////////////////////////////////////////////// output of im_X1_15

q[271]= (im_X11_0 * p_cos_0 );
q[272]= (im_X12_0 * p_cos_216 );
q[273]= (im_X13_0 * p_cos_72 );
q[274]= (im_X14_0 * p_cos_288 );
q[275]= (im_X15_0 * p_cos_144 );
q[276]= (re_X12_0 * p_sin_216 );
q[277]= (re_X13_0 * p_sin_72 );
q[278]= (re_X14_0 * p_sin_288 );
q[279]= (re_X15_0 * p_sin_144 );

p[270] = q[270][31:16] + q[270][15];
p[271] = q[271][31:16] + q[271][15];
p[272] = q[272][31:16] + q[272][15];
p[273] = q[273][31:16] + q[273][15];
p[274] = q[274][31:16] + q[274][15];
p[275] = q[275][31:16] + q[275][15];
p[276] = q[276][31:16] + q[276][15];
p[277] = q[277][31:16] + q[277][15];
p[278] = q[278][31:16] + q[278][15];
p[279] = q[279][31:16] + q[279][15];

/////////////////////////////////////////////////////////////////////////////////// output of re_X1_16

q[280]= (re_X11_1 * p_cos_0 );
q[281]= (re_X12_1 * p_cos_230_4 );
q[282]= (re_X13_1 * p_cos_100_8 );
q[283]= (re_X14_1 * p_cos_331_2 );
q[284]= (re_X15_1 * p_cos_201_6 );
q[285]= (im_X12_1 * p_sin_230_4 );
q[286]= (im_X13_1 * p_sin_100_8 );
q[287]= (im_X14_1 * p_sin_331_2 );
q[288]= (im_X15_1 * p_sin_201_6 );

p[280] = q[280][31:16] + q[280][15];
p[281] = q[281][31:16] + q[281][15];
p[282] = q[282][31:16] + q[282][15];
p[283] = q[283][31:16] + q[283][15];
p[284] = q[284][31:16] + q[284][15];
p[285] = q[285][31:16] + q[285][15];
p[286] = q[286][31:16] + q[286][15];
p[287] = q[287][31:16] + q[287][15];
p[288] = q[288][31:16] + q[288][15];


////////////////////////////////////////////////////////////////////////////////// output of im_X1_16

q[289]= (im_X11_1 * p_cos_0 );
q[290]= (im_X12_1 * p_cos_230_4 );
q[291]= (im_X13_1 * p_cos_100_8 );
q[292]= (im_X14_1 * p_cos_331_2 );
q[293]= (im_X15_1 * p_cos_201_6 );
q[294]= (re_X12_1 * p_sin_230_4 );
q[295]= (re_X13_1 * p_sin_100_8 );
q[296]= (re_X14_1 * p_sin_331_2 );
q[297]= (re_X15_1 * p_sin_201_6 );

p[289] = q[289][31:16] + q[289][15];
p[290] = q[290][31:16] + q[290][15];
p[291] = q[291][31:16] + q[291][15];
p[292] = q[292][31:16] + q[292][15];
p[293] = q[293][31:16] + q[293][15];
p[294] = q[294][31:16] + q[294][15];
p[295] = q[295][31:16] + q[295][15];
p[296] = q[296][31:16] + q[296][15];
p[297] = q[297][31:16] + q[297][15];

////////////////////////////////////////////////////////////////////////////////// output of re_X1_17

q[298]= (re_X11_2 * p_cos_0 );
q[299]= (re_X12_2 * p_cos_244_8 );
q[300]= (re_X13_2 * p_cos_129_6 );
q[301]= (re_X14_2 * p_cos_14_4 );
q[302]= (re_X15_2 * p_cos_259_2 );
q[303]= (im_X12_2 * p_sin_244_8 );
q[304]= (im_X13_2 * p_sin_129_6 );
q[305]= (im_X14_2 * p_sin_14_4 );
q[306]= (im_X15_2 * p_sin_259_2 );

p[298] = q[298][31:16] + q[298][15];
p[299] = q[299][31:16] + q[299][15];
p[300] = q[300][31:16] + q[300][15];
p[301] = q[301][31:16] + q[301][15];
p[302] = q[302][31:16] + q[302][15];
p[303] = q[303][31:16] + q[303][15];
p[304] = q[304][31:16] + q[304][15];
p[305] = q[305][31:16] + q[305][15];
p[306] = q[306][31:16] + q[306][15];

/////////////////////////////////////////////////////////////////////////////////// output of im_X1_17

q[307]= (im_X11_2 * p_cos_0 );
q[308]= (im_X12_2 * p_cos_244_8 );
q[309]= (im_X13_2 * p_cos_129_6 );
q[310]= (im_X14_2 * p_cos_14_4 );
q[311]= (im_X15_2 * p_cos_259_2 );
q[312]= (re_X12_2 * p_sin_244_8 );
q[313]= (re_X13_2 * p_sin_129_6 );
q[314]= (re_X14_2 * p_sin_14_4 );
q[315]= (re_X15_2 * p_sin_259_2 );

p[307] = q[307][31:16] + q[307][15];
p[308] = q[308][31:16] + q[308][15];
p[309] = q[309][31:16] + q[309][15];
p[310] = q[310][31:16] + q[310][15];
p[311] = q[311][31:16] + q[311][15];
p[312] = q[312][31:16] + q[312][15];
p[313] = q[313][31:16] + q[313][15];
p[314] = q[314][31:16] + q[314][15];
p[315] = q[315][31:16] + q[315][15];

////////////////////////////////////////////////////////////////////////////////// output of re_X1_18

q[316]= (re_X11_3 * p_cos_0 );
q[317]= (re_X12_3 * p_cos_259_2 );
q[318]= (re_X13_3 * p_cos_158_4 );
q[319]= (re_X14_3 * p_cos_57_6 );
q[320]= (re_X15_3 * p_cos_316_8 );
q[321]= (im_X12_3 * p_sin_259_2 );
q[322]= (im_X13_3 * p_sin_158_4 );
q[323]= (im_X14_3 * p_sin_57_6 );
q[324]= (im_X15_3 * p_sin_316_8 );

p[316] = q[316][31:16] + q[316][15];
p[317] = q[317][31:16] + q[317][15];
p[318] = q[318][31:16] + q[318][15];
p[319] = q[319][31:16] + q[319][15];
p[320] = q[320][31:16] + q[320][15];
p[321] = q[321][31:16] + q[321][15];
p[322] = q[322][31:16] + q[322][15];
p[323] = q[323][31:16] + q[323][15];
p[324] = q[324][31:16] + q[324][15];

/////////////////////////////////////////////////////////////////////////////// output of im_X1_18

q[325]= (im_X11_3 * p_cos_0 );
q[326]= (im_X12_3 * p_cos_259_2 );
q[327]= (im_X13_3 * p_cos_158_4 );
q[328]= (im_X14_3 * p_cos_57_6 );
q[329]= (im_X15_3 * p_cos_316_8 );
q[330]= (re_X12_3 * p_sin_259_2 );
q[331]= (re_X13_3 * p_sin_158_4 );
q[332]= (re_X14_3 * p_sin_57_6 );
q[333]= (re_X15_3 * p_sin_316_8 );

p[325] = q[325][31:16] + q[325][15];
p[326] = q[326][31:16] + q[326][15];
p[327] = q[327][31:16] + q[327][15];
p[328] = q[328][31:16] + q[328][15];
p[329] = q[329][31:16] + q[329][15];
p[330] = q[330][31:16] + q[330][15];
p[331] = q[331][31:16] + q[331][15];
p[332] = q[332][31:16] + q[332][15];
p[333] = q[333][31:16] + q[333][15];

/////////////////////////////////////////////////////////////////////////////// output of re_X1_19

q[334]= (re_X11_4 * p_cos_0 );
q[335]= (re_X12_4 * p_cos_273_6 );
q[336]= (re_X13_4 * p_cos_187_2 );
q[337]= (re_X14_4 * p_cos_100_8 );
q[338]= (re_X15_4 * p_cos_14_4 );
q[339]= (im_X12_4 * p_sin_273_6 );
q[340]= (im_X13_4 * p_sin_187_2 );
q[341]= (im_X14_4 * p_sin_100_8 );
q[342]= (im_X15_4 * p_sin_14_4 );

p[334] = q[334][31:16] + q[334][15];
p[335] = q[335][31:16] + q[335][15];
p[336] = q[336][31:16] + q[336][15];
p[337] = q[337][31:16] + q[337][15];
p[338] = q[338][31:16] + q[338][15];
p[339] = q[339][31:16] + q[339][15];
p[340] = q[340][31:16] + q[340][15];
p[341] = q[341][31:16] + q[341][15];
p[342] = q[342][31:16] + q[342][15];

/////////////////////////////////////////////////////////////////////////////// output of im_X1_19

q[343]= (im_X11_4 * p_cos_0 );
q[344]= (im_X12_4 * p_cos_273_6 );
q[345]= (im_X13_4 * p_cos_187_2 );
q[346]= (im_X14_4 * p_cos_100_8 );
q[347]= (im_X15_4 * p_cos_14_4 );
q[348]= (re_X12_4 * p_sin_273_6 );
q[349]= (re_X13_4 * p_sin_187_2 );
q[350]= (re_X14_4 * p_sin_100_8 );
q[351]= (re_X15_4 * p_sin_14_4 );

p[343] = q[343][31:16] + q[343][15];
p[344] = q[344][31:16] + q[344][15];
p[345] = q[345][31:16] + q[345][15];
p[346] = q[346][31:16] + q[346][15];
p[347] = q[347][31:16] + q[347][15];
p[348] = q[348][31:16] + q[348][15];
p[349] = q[349][31:16] + q[349][15];
p[350] = q[350][31:16] + q[350][15];
p[351] = q[351][31:16] + q[351][15];

////////////////////////////////////////////////////////////////////////////// output of re_X1_20

q[352]= (re_X11_0 * p_cos_0 );
q[353]= (re_X12_0 * p_cos_288 );
q[354]= (re_X13_0 * p_cos_216 );
q[355]= (re_X14_0 * p_cos_144 );
q[356]= (re_X15_0 * p_cos_72 );
q[357]= (im_X12_0 * p_sin_288 );
q[358]= (im_X13_0 * p_sin_216);
q[359]= (im_X14_0 * p_sin_144 );
q[360]= (im_X15_0 * p_sin_72 );

p[352] = q[352][31:16] + q[352][15];
p[353] = q[353][31:16] + q[353][15];
p[354] = q[354][31:16] + q[354][15];
p[355] = q[355][31:16] + q[355][15];
p[356] = q[356][31:16] + q[356][15];
p[357] = q[357][31:16] + q[357][15];
p[358] = q[358][31:16] + q[358][15];
p[359] = q[359][31:16] + q[359][15];
p[360] = q[360][31:16] + q[360][15];

/////////////////////////////////////////////////////////////////////////////// output of im_X1_20

q[361]= (im_X11_0 * p_cos_0 );
q[362]= (im_X12_0 * p_cos_288 );
q[363]= (im_X13_0 * p_cos_216 );
q[364]= (im_X14_0 * p_cos_144 );
q[365]= (im_X15_0 * p_cos_72 );
q[366]= (re_X12_0 * p_sin_288 );
q[367]= (re_X13_0 * p_sin_216 );
q[368]= (re_X14_0 * p_sin_144 );
q[369]= (re_X15_0 * p_sin_72 );

p[361] = q[361][31:16] + q[361][15];
p[362] = q[362][31:16] + q[362][15];
p[363] = q[363][31:16] + q[363][15];
p[364] = q[364][31:16] + q[364][15];
p[365] = q[365][31:16] + q[365][15];
p[366] = q[366][31:16] + q[366][15];
p[367] = q[367][31:16] + q[367][15];
p[368] = q[368][31:16] + q[368][15];
p[369] = q[369][31:16] + q[369][15];

/////////////////////////////////////////////////////////////////////////////// output of re_X1_21

q[370]= (re_X11_1 * p_cos_0 );
q[371]= (re_X12_1 * p_cos_302_4 );
q[372]= (re_X13_1 * p_cos_244_8 );
q[373]= (re_X14_1 * p_cos_187_2 );
q[374]= (re_X15_1 * p_cos_129_6 );
q[375]= (im_X12_1 * p_sin_302_4 );
q[376]= (im_X13_1 * p_sin_244_8 );
q[377]= (im_X14_1 * p_sin_187_2 );
q[378]= (im_X15_1 * p_sin_129_6 );

p[370] = q[370][31:16] + q[370][15];
p[371] = q[371][31:16] + q[371][15];
p[372] = q[372][31:16] + q[372][15];
p[373] = q[373][31:16] + q[373][15];
p[374] = q[374][31:16] + q[374][15];
p[375] = q[375][31:16] + q[375][15];
p[376] = q[376][31:16] + q[376][15];
p[377] = q[377][31:16] + q[377][15];
p[378] = q[378][31:16] + q[378][15];

/////////////////////////////////////////////////////////////////////////////// output of im_X1_21

q[379]= (im_X11_1 * p_cos_0 );
q[380]= (im_X12_1 * p_cos_302_4 );
q[381]= (im_X13_1 * p_cos_244_8 );
q[382]= (im_X14_1 * p_cos_187_2 );
q[383]= (im_X15_1 * p_cos_129_6 );
q[384]= (re_X12_1 * p_sin_302_4 );
q[385]= (re_X13_1 * p_sin_244_8 );
q[386]= (re_X14_1 * p_sin_187_2 );
q[387]= (re_X15_1 * p_sin_129_6 );

p[379] = q[379][31:16] + q[379][15];
p[380] = q[380][31:16] + q[380][15];
p[381] = q[381][31:16] + q[381][15];
p[382] = q[382][31:16] + q[382][15];
p[383] = q[383][31:16] + q[383][15];
p[384] = q[384][31:16] + q[384][15];
p[385] = q[385][31:16] + q[385][15];
p[386] = q[386][31:16] + q[386][15];
p[387] = q[387][31:16] + q[387][15];

/////////////////////////////////////////////////////////////////////////////// output of re_X1_22

q[388]= (re_X11_2 * p_cos_0 );
q[389]= (re_X12_2 * p_cos_316_8 );
q[390]= (re_X13_2 * p_cos_273_6 );
q[391]= (re_X14_2 * p_cos_230_4 );
q[392]= (re_X15_2 * p_cos_187_2 );
q[393]= (im_X12_2 * p_sin_316_8 );
q[394]= (im_X13_2 * p_sin_273_6 );
q[395]= (im_X14_2 * p_sin_230_4 );
q[396]= (im_X15_2 * p_sin_187_2 );

p[388] = q[388][31:16] + q[388][15];
p[389] = q[389][31:16] + q[389][15];
p[390] = q[390][31:16] + q[390][15];
p[391] = q[391][31:16] + q[391][15];
p[392] = q[392][31:16] + q[392][15];
p[393] = q[393][31:16] + q[393][15];
p[394] = q[394][31:16] + q[394][15];
p[395] = q[395][31:16] + q[395][15];
p[396] = q[396][31:16] + q[396][15];

/////////////////////////////////////////////////////////////////////////////// output of im_X1_22

q[397]= (im_X11_2 * p_cos_0 );
q[398]= (im_X12_2 * p_cos_316_8 );
q[399]= (im_X13_2 * p_cos_273_6 );
q[400]= (im_X14_2 * p_cos_230_4 );
q[401]= (im_X15_2 * p_cos_187_2 );
q[402]= (re_X12_2 * p_sin_316_8 );
q[403]= (re_X13_2 * p_sin_273_6 );
q[404]= (re_X14_2 * p_sin_230_4 );
q[405]= (re_X15_2 * p_sin_187_2 );

p[397] = q[397][31:16] + q[397][15];
p[398] = q[398][31:16] + q[398][15];
p[399] = q[399][31:16] + q[399][15];
p[400] = q[400][31:16] + q[400][15];
p[401] = q[401][31:16] + q[401][15];
p[402] = q[402][31:16] + q[402][15];
p[403] = q[403][31:16] + q[403][15];
p[404] = q[404][31:16] + q[404][15];
p[405] = q[405][31:16] + q[405][15];

//////////////////////////////////////////////////////////////////////////////// output of re_X1_23

q[406]= (re_X11_3 * p_cos_0 );
q[407]= (re_X12_3 * p_cos_331_2 );
q[408]= (re_X13_3 * p_cos_302_4 );
q[409]= (re_X14_3 * p_cos_273_6 );
q[410]= (re_X15_3 * p_cos_244_8 );
q[411]= (im_X12_3 * p_sin_331_2 );
q[412]= (im_X13_3 * p_sin_302_4 );
q[413]= (im_X14_3 * p_sin_273_6 );
q[414]= (im_X15_3 * p_sin_244_8 );

p[406] = q[406][31:16] + q[406][15];
p[407] = q[407][31:16] + q[407][15];
p[408] = q[408][31:16] + q[408][15];
p[409] = q[409][31:16] + q[409][15];
p[410] = q[410][31:16] + q[410][15];
p[411] = q[411][31:16] + q[411][15];
p[412] = q[412][31:16] + q[412][15];
p[413] = q[413][31:16] + q[413][15];
p[414] = q[414][31:16] + q[414][15];

//////////////////////////////////////////////////////////////////////////////// output of im_X1_23

q[415]= (im_X11_3 * p_cos_0 );
q[416]= (im_X12_3 * p_cos_331_2 );
q[417]= (im_X13_3 * p_cos_302_4 );
q[418]= (im_X14_3 * p_cos_273_6 );
q[419]= (im_X15_3 * p_cos_244_8 );
q[420]= (re_X12_3 * p_sin_331_2 );
q[421]= (re_X13_3 * p_sin_302_4 );
q[422]= (re_X14_3 * p_sin_273_6 );
q[423]= (re_X15_3 * p_sin_244_8 );

p[415] = q[415][31:16] + q[415][15];
p[416] = q[416][31:16] + q[416][15];
p[417] = q[417][31:16] + q[417][15];
p[418] = q[418][31:16] + q[418][15];
p[419] = q[419][31:16] + q[419][15];
p[420] = q[420][31:16] + q[420][15];
p[421] = q[421][31:16] + q[421][15];
p[422] = q[422][31:16] + q[422][15];
p[423] = q[423][31:16] + q[423][15];

///////////////////////////////////////////////////////////////////////////////// output of re_X1_24

q[424]= (re_X11_4 * p_cos_0 );
q[425]= (re_X12_4 * p_cos_345_6 );
q[426]= (re_X13_4 * p_cos_331_2 );
q[427]= (re_X14_4 * p_cos_316_8 );
q[428]= (re_X15_4 * p_cos_302_4 );
q[429]= (im_X12_4 * p_sin_345_6 );
q[430]= (im_X13_4 * p_sin_331_2 );
q[431]= (im_X14_4 * p_sin_316_8 );
q[432]= (im_X15_4 * p_sin_302_4 );

p[424] = q[424][31:16] + q[424][15];
p[425] = q[425][31:16] + q[425][15];
p[426] = q[426][31:16] + q[426][15];
p[427] = q[427][31:16] + q[427][15];
p[428] = q[428][31:16] + q[428][15];
p[429] = q[429][31:16] + q[429][15];
p[430] = q[430][31:16] + q[430][15];
p[431] = q[431][31:16] + q[431][15];
p[432] = q[432][31:16] + q[432][15];

///////////////////////////////////////////////////////////////////////////////// output of im_X1_24

q[433]= (im_X11_4 * p_cos_0 );
q[434]= (im_X12_4 * p_cos_345_6 );
q[435]= (im_X13_4 * p_cos_331_2 );
q[436]= (im_X14_4 * p_cos_316_8 );
q[437]= (im_X15_4 * p_cos_302_4 );
q[438]= (re_X12_4 * p_sin_345_6 );
q[439]= (re_X13_4 * p_sin_331_2 );
q[440]= (re_X14_4 * p_sin_316_8 );
q[441]= (re_X15_4 * p_sin_302_4 );

p[433] = q[433][31:16] + q[433][15];
p[434] = q[434][31:16] + q[434][15];
p[435] = q[435][31:16] + q[435][15];
p[436] = q[436][31:16] + q[436][15];
p[437] = q[437][31:16] + q[437][15];
p[438] = q[438][31:16] + q[438][15];
p[439] = q[439][31:16] + q[439][15];
p[440] = q[440][31:16] + q[440][15];
p[441] = q[441][31:16] + q[441][15];



m[0] = div_5*(p[0] + p[1] + p[2] + p[3] + p[4]);
m[1] = div_5*(p[5] + p[6] + p[7] + p[8] + p[9]);
m[2] = div_5*(p[10] + p[11] + p[12] + p[13] + p[14] + p[15] + p[16] + p[17] + p[18]);
m[3] = div_5*(p[19] + p[20] + p[21] + p[22] + p[23] - p[24] - p[25] - p[26] - p[27]);
m[4] = div_5*(p[28] + p[29] + p[30] + p[31] + p[32] + p[33] + p[34] + p[35] + p[36]);
m[5] = div_5*(p[37] + p[38] + p[39] + p[40] + p[41] - p[42] - p[43] - p[44] - p[45]);
m[6] = div_5*(p[46] + p[47] + p[48] + p[49] + p[50] + p[51] + p[52] + p[53] + p[54]);
m[7] = div_5*(p[55] + p[56] + p[57] + p[58] + p[59] - p[60] - p[61] - p[62] - p[63]);
m[8] = div_5*(p[64] + p[65] + p[66] + p[67] + p[68] + p[69] + p[70] + p[71] + p[72]);
m[9] = div_5*(p[73] + p[74] + p[75] + p[76] + p[77] - p[78] - p[79] - p[80] - p[81]);
m[10] = div_5*(p[82] + p[83] + p[84] + p[85] + p[86] + p[87] + p[88] + p[89] + p[90]);
m[11] = div_5*(p[91] + p[92] + p[93] + p[94] + p[95] - p[96] - p[97] - p[98] - p[99]);
m[12] = div_5*(p[100] + p[101] + p[102] + p[103] + p[104] + p[105] + p[106] + p[107] + p[108]);
m[13] = div_5*(p[109] + p[110] + p[111] + p[112] + p[113] - p[114] - p[115] - p[116] - p[117]);
m[14] = div_5*(p[118] + p[119] + p[120] + p[121] + p[122] + p[123] + p[124] + p[125] + p[126]);
m[15] = div_5*(p[127] + p[128] + p[129] + p[130] + p[131] - p[132] - p[133] - p[134] - p[135]);
m[16] = div_5*(p[136] + p[137] + p[138] + p[139] + p[140] + p[141] + p[142] + p[143] + p[144]);
m[17] = div_5*(p[145] + p[146] + p[147] + p[148] + p[149] - p[150] - p[151] - p[152] - p[153]);
m[18] = div_5*(p[154] + p[155] + p[156] + p[157] + p[158] + p[159] + p[160] + p[161] + p[162]);
m[19] = div_5*(p[163] + p[164] + p[165] + p[166] + p[167] - p[168] - p[169] - p[170] - p[171]);
m[20] = div_5*(p[172] + p[173] + p[174] + p[175] + p[176] + p[177] + p[178] + p[179] + p[180]);
m[21] = div_5*(p[181] + p[182] + p[183] + p[184] + p[185] - p[186] - p[187] - p[188] - p[189]);
m[22]= div_5*(p[190] + p[191] + p[192] + p[193] + p[194] + p[195] + p[196] + p[197] + p[198]);
m[23]= div_5*(p[199] + p[200] + p[201] + p[202] + p[203] - p[204] - p[205] - p[206] - p[207]);
m[24]= div_5*(p[208] + p[209] + p[210] + p[211] + p[212] + p[213] + p[214] + p[215] + p[216]);
m[25]= div_5*(p[217] + p[218] + p[219] + p[220] + p[221] - p[222] - p[223] - p[224] - p[225]);
m[26]= div_5*(p[226] + p[227] + p[228] + p[229] + p[230] + p[231] + p[232] + p[233] + p[234]);
m[27]= div_5*(p[235] + p[236] + p[237] + p[238] + p[239] - p[240] - p[241] - p[242] - p[243]);
m[28]= div_5*(p[244] + p[245] + p[246] + p[247] + p[248] + p[249] + p[250] + p[251] + p[252]);
m[29]= div_5*(p[253] + p[254] + p[255] + p[256] + p[257] - p[258] - p[259] - p[260] - p[261]);
m[30]= div_5*(p[262] + p[263] + p[264] + p[265] + p[266] + p[267] + p[268] + p[269] + p[270]);
m[31]= div_5*(p[271] + p[272] + p[273] + p[274] + p[275] - p[276] - p[277] - p[278] - p[279]);
m[32]= div_5*(p[280] + p[281] + p[282] + p[283] + p[284] + p[285] + p[286] + p[287] + p[288]);
m[33]= div_5*(p[289] + p[290] + p[291] + p[292] + p[293] - p[294] - p[295] - p[296] - p[297]);
m[34]= div_5*(p[298] + p[299] + p[300] + p[301] + p[302] + p[303] + p[304] + p[305] + p[306]);
m[35]= div_5*(p[307] + p[308] + p[309] + p[310] + p[311] - p[312] - p[313] - p[314] - p[315]);
m[36]= div_5*(p[316] + p[317] + p[318] + p[319] + p[320] + p[321] + p[322] + p[323] + p[324]);
m[37]= div_5*(p[325] + p[326] + p[327] + p[328] + p[329] - p[330] - p[331] - p[332] - p[333]);
m[38]= div_5*(p[334] + p[335] + p[336] + p[337] + p[338] + p[339] + p[340] + p[341] + p[342]);
m[39]= div_5*(p[343] + p[344] + p[345] + p[346] + p[347] - p[348] - p[349] - p[350] - p[351]);
m[40]= div_5*(p[352] + p[353] + p[354] + p[355] + p[356] + p[357] + p[358] + p[359] + p[360]);
m[41]= div_5*(p[361] + p[362] + p[363] + p[364] + p[365] - p[366] - p[367] - p[368] - p[369]);
m[42]= div_5*(p[370] + p[371] + p[372] + p[373] + p[374] + p[375] + p[376] + p[377] + p[378]);
m[43]= div_5*(p[379] + p[380] + p[381] + p[382] + p[383] - p[384] - p[385] - p[386] - p[387]);
m[44]= div_5*(p[388] + p[389] + p[390] + p[391] + p[392] + p[393] + p[394] + p[395] + p[396]);
m[45]= div_5*(p[397] + p[398] + p[399] + p[400] + p[401] - p[402] - p[403] - p[404] - p[405]);
m[46]= div_5*(p[406] + p[407] + p[408] + p[409] + p[410] + p[411] + p[412] + p[413] + p[414]);
m[47]= div_5*(p[415] + p[416] + p[417] + p[418] + p[419] - p[420] - p[421] - p[422] - p[423]);
m[48]= div_5*(p[424] + p[425] + p[426] + p[427] + p[428] + p[429] + p[430] + p[431] + p[432]);
m[49]= div_5*(p[433] + p[434] + p[435] + p[436] + p[437] - p[438] - p[439] - p[440] - p[441]);


re_X1_0 = m[0][28:12] + m[0][11];
im_X1_0 = m[1][28:12] + m[1][11];
re_X1_1 = m[2][28:12] + m[2][11] ;
 im_X1_1 = m[3][28:12] + m[3][11];
re_X1_2 = m[4][28:12] + m[4][11] ;
 im_X1_2 = m[5][28:12] + m[5][11];
re_X1_3 = m[6][28:12] + m[6][11] ;
 im_X1_3 = m[7][28:12] + m[7][11];
re_X1_4 = m[8][28:12] + m[8][11] ;
 im_X1_4 = m[9][28:12] + m[9][11];
re_X1_5 = m[10][28:12] + m[10][11] ;
 im_X1_5 = m[11][28:12] + m[11][11];
re_X1_6 = m[12][28:12] + m[12][11] ;
 im_X1_6 = m[13][28:12] + m[13][11];
re_X1_7 = m[14][28:12] + m[14][11] ;
 im_X1_7 = m[15][28:12] + m[15][11];
re_X1_8 = m[16][28:12] + m[16][11] ;
 im_X1_8 = m[17][28:12] + m[17][11];
re_X1_9 = m[18][28:12] + m[18][11] ;
 im_X1_9 = m[19][28:12] + m[19][11];
re_X1_10 = m[20][28:12] + m[20][11] ;
 im_X1_10 = m[21][28:12] + m[21][11];
re_X1_11 = m[22][28:12] + m[22][11] ;
 im_X1_11 = m[23][28:12] + m[23][11];
re_X1_12 = m[24][28:12] + m[24][11] ;
 im_X1_12 = m[25][28:12] + m[25][11];
re_X1_13 = m[26][28:12] + m[26][11] ;
 im_X1_13 = m[27][28:12] + m[27][11];
re_X1_14 = m[28][28:12] + m[28][11] ;
 im_X1_14 = m[29][28:12] + m[29][11];
re_X1_15 = m[30][28:12] + m[30][11] ;
 im_X1_15 = m[31][28:12] + m[31][11];
re_X1_16 = m[32][28:12] + m[32][11] ;
 im_X1_16 = m[33][28:12] + m[33][11];
re_X1_17 = m[34][28:12] + m[34][11] ;
 im_X1_17 = m[35][28:12] + m[35][11];
re_X1_18 = m[36][28:12] + m[36][11] ;
 im_X1_18 = m[37][28:12] + m[37][11];
re_X1_19 = m[38][28:12] + m[38][11] ;
 im_X1_19 = m[39][28:12] + m[39][11];
re_X1_20 = m[40][28:12] + m[40][11] ;
 im_X1_20 = m[41][28:12] + m[41][11];
re_X1_21 = m[42][28:12] + m[42][11] ;
 im_X1_21 = m[43][28:12] + m[43][11];
re_X1_22 = m[44][28:12] + m[44][11] ;
 im_X1_22 = m[45][28:12] + m[45][11];
re_X1_23 = m[46][28:12] + m[46][11] ;
 im_X1_23 = m[47][28:12] + m[47][11];
re_X1_24 = m[48][28:12] + m[48][11] ;
 im_X1_24 = m[49][28:12] + m[49][11];
end

endmodule

////////////////FINAL FFT MODULE////////////////////

module FFT(clk,re_x_0,im_x_0,re_x_1,im_x_1,re_x_2,im_x_2,re_x_3,im_x_3,re_x_4,im_x_4,re_x_5,im_x_5,re_x_6,im_x_6,re_x_7,im_x_7,re_x_8,im_x_8,re_x_9,im_x_9,re_x_10,im_x_10,
re_x_11,im_x_11,re_x_12,im_x_12,re_x_13,im_x_13,re_x_14,im_x_14,re_x_15,im_x_15,re_x_16,im_x_16,re_x_17,im_x_17,re_x_18,im_x_18,re_x_19,im_x_19,re_x_20,im_x_20,
re_x_21,im_x_21,re_x_22,im_x_22,re_x_23,im_x_23,re_x_24,im_x_24,re_x_25,im_x_25,re_x_26,im_x_26,re_x_27,im_x_27,re_x_28,im_x_28,re_x_29,im_x_29,re_x_30,im_x_30,
re_x_31,im_x_31,re_x_32,im_x_32,re_x_33,im_x_33,re_x_34,im_x_34,re_x_35,im_x_35,re_x_36,im_x_36,re_x_37,im_x_37,re_x_38,im_x_38,re_x_39,im_x_39,re_x_40,im_x_40,
re_x_41,im_x_41,re_x_42,im_x_42,re_x_43,im_x_43,re_x_44,im_x_44,re_x_45,im_x_45,re_x_46,im_x_46,re_x_47,im_x_47,re_x_48,im_x_48,re_x_49,im_x_49,
re_X_0,im_X_0,re_X_1,im_X_1,re_X_2,im_X_2,re_X_3,im_X_3,re_X_4,im_X_4,re_X_5,im_X_5,re_X_6,im_X_6,re_X_7,im_X_7,re_X_8,im_X_8,re_X_9,im_X_9,re_X_10,im_X_10,
re_X_11,im_X_11,re_X_12,im_X_12,re_X_13,im_X_13,re_X_14,im_X_14,re_X_15,im_X_15,re_X_16,im_X_16,re_X_17,im_X_17,re_X_18,im_X_18,re_X_19,im_X_19,re_X_20,im_X_20,
re_X_21,im_X_21,re_X_22,im_X_22,re_X_23,im_X_23,re_X_24,im_X_24,re_X_25,im_X_25,re_X_26,im_X_26,re_X_27,im_X_27,re_X_28,im_X_28,re_X_29,im_X_29,re_X_30,im_X_30,
re_X_31,im_X_31,re_X_32,im_X_32,re_X_33,im_X_33,re_X_34,im_X_34,re_X_35,im_X_35,re_X_36,im_X_36,re_X_37,im_X_37,re_X_38,im_X_38,re_X_39,im_X_39,re_X_40,im_X_40,
re_X_41,im_X_41,re_X_42,im_X_42,re_X_43,im_X_43,re_X_44,im_X_44,re_X_45,im_X_45,re_X_46,im_X_46,re_X_47,im_X_47,re_X_48,im_X_48,re_X_49,im_X_49);

input signed [15:0] re_x_0,im_x_0,re_x_1,im_x_1,re_x_2,im_x_2,re_x_3,im_x_3,re_x_4,im_x_4,re_x_5,im_x_5,re_x_6,im_x_6,re_x_7,im_x_7,re_x_8,im_x_8,re_x_9,im_x_9,re_x_10,im_x_10,
re_x_11,im_x_11,re_x_12,im_x_12,re_x_13,im_x_13,re_x_14,im_x_14,re_x_15,im_x_15,re_x_16,im_x_16,re_x_17,im_x_17,re_x_18,im_x_18,re_x_19,im_x_19,re_x_20,im_x_20,
re_x_21,im_x_21,re_x_22,im_x_22,re_x_23,im_x_23,re_x_24,im_x_24,re_x_25,im_x_25,re_x_26,im_x_26,re_x_27,im_x_27,re_x_28,im_x_28,re_x_29,im_x_29,re_x_30,im_x_30,
re_x_31,im_x_31,re_x_32,im_x_32,re_x_33,im_x_33,re_x_34,im_x_34,re_x_35,im_x_35,re_x_36,im_x_36,re_x_37,im_x_37,re_x_38,im_x_38,re_x_39,im_x_39,re_x_40,im_x_40,
re_x_41,im_x_41,re_x_42,im_x_42,re_x_43,im_x_43,re_x_44,im_x_44,re_x_45,im_x_45,re_x_46,im_x_46,re_x_47,im_x_47,re_x_48,im_x_48,re_x_49,im_x_49;

input clk;

output signed [15:0] re_X_0,im_X_0,re_X_1,im_X_1,re_X_2,im_X_2,re_X_3,im_X_3,re_X_4,im_X_4,re_X_5,im_X_5,re_X_6,im_X_6,re_X_7,im_X_7,re_X_8,im_X_8,re_X_9,im_X_9,re_X_10,im_X_10,
re_X_11,im_X_11,re_X_12,im_X_12,re_X_13,im_X_13,re_X_14,im_X_14,re_X_15,im_X_15,re_X_16,im_X_16,re_X_17,im_X_17,re_X_18,im_X_18,re_X_19,im_X_19,re_X_20,im_X_20,
re_X_21,im_X_21,re_X_22,im_X_22,re_X_23,im_X_23,re_X_24,im_X_24,re_X_25,im_X_25,re_X_26,im_X_26,re_X_27,im_X_27,re_X_28,im_X_28,re_X_29,im_X_29,re_X_30,im_X_30,
re_X_31,im_X_31,re_X_32,im_X_32,re_X_33,im_X_33,re_X_34,im_X_34,re_X_35,im_X_35,re_X_36,im_X_36,re_X_37,im_X_37,re_X_38,im_X_38,re_X_39,im_X_39,re_X_40,im_X_40,
re_X_41,im_X_41,re_X_42,im_X_42,re_X_43,im_X_43,re_X_44,im_X_44,re_X_45,im_X_45,re_X_46,im_X_46,re_X_47,im_X_47,re_X_48,im_X_48,re_X_49,im_X_49;

real re_X2_2_fractional,im_X2_2_fractional,re_X1_2_fractional,re_X21_2_fractional,re_X22_2_fractional,re_X23_2_fractional,re_X24_2_fractional,re_X25_2_fractional,im_X21_2_fractional,
im_X22_2_fractional,im_X23_2_fractional,im_X24_2_fractional,im_X25_2_fractional;

wire signed [16:0] re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4,re_X12_0,im_X12_0,re_X12_1,im_X12_1,re_X12_2,im_X12_2,re_X12_3,im_X12_3,re_X12_4,
im_X12_4,re_X13_0,im_X13_0,re_X13_1,im_X13_1,re_X13_2,im_X13_2,re_X13_3,im_X13_3,re_X13_4,im_X13_4,re_X14_0,im_X14_0,re_X14_1,im_X14_1,re_X14_2,im_X14_2,re_X14_3,im_X14_3,re_X14_4,im_X14_4,
re_X15_0,im_X15_0,re_X15_1,im_X15_1,re_X15_2,im_X15_2,re_X15_3,im_X15_3,re_X15_4,im_X15_4,re_X21_0,im_X21_0,re_X21_1,im_X21_1,re_X21_2,im_X21_2,re_X21_3,im_X21_3,re_X21_4,im_X21_4,
re_X22_0,im_X22_0,re_X22_1,im_X22_1,re_X22_2,im_X22_2,re_X22_3,im_X22_3,re_X22_4,im_X22_4,re_X23_0,im_X23_0,re_X23_1,im_X23_1,re_X23_2,im_X23_2,re_X23_3,im_X23_3,re_X23_4,im_X23_4,
re_X24_0,im_X24_0,re_X24_1,im_X24_1,re_X24_2,im_X24_2,re_X24_3,im_X24_3,re_X24_4,im_X24_4,re_X25_0,im_X25_0,re_X25_1,im_X25_1,re_X25_2,im_X25_2,re_X25_3,im_X25_3,re_X25_4,im_X25_4;

wire signed [16:0] re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,
im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,
re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24,re_X2_0,im_X2_0,re_X2_1,im_X2_1,re_X2_2,im_X2_2,re_X2_3,im_X2_3,re_X2_4,im_X2_4,
re_X2_5,im_X2_5,re_X2_6,im_X2_6,re_X2_7,im_X2_7,re_X2_8,im_X2_8,re_X2_9,im_X2_9,re_X2_10,im_X2_10,re_X2_11,im_X2_11,re_X2_12,im_X2_12,re_X2_13,im_X2_13,re_X2_14,im_X2_14,re_X2_15,im_X2_15,
re_X2_16,im_X2_16,re_X2_17,im_X2_17,re_X2_18,im_X2_18,re_X2_19,im_X2_19,re_X2_20,im_X2_20,re_X2_21,im_X2_21,re_X2_22,im_X2_22,re_X2_23,im_X2_23,re_X2_24,im_X2_24;


///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


fft_radix5 FFT1(clk,re_x_0,re_x_10,re_x_20,re_x_30,re_x_40,im_x_0,im_x_10,im_x_20,im_x_30,im_x_40,re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4);
fft_radix5 FFT2(clk,re_x_2,re_x_12,re_x_22,re_x_32,re_x_42,im_x_2,im_x_12,im_x_22,im_x_32,im_x_42,re_X12_0,im_X12_0,re_X12_1,im_X12_1,re_X12_2,im_X12_2,re_X12_3,im_X12_3,re_X12_4,im_X12_4);
fft_radix5 FFT3(clk,re_x_4,re_x_14,re_x_24,re_x_34,re_x_44,im_x_4,im_x_14,im_x_24,im_x_34,im_x_44,re_X13_0,im_X13_0,re_X13_1,im_X13_1,re_X13_2,im_X13_2,re_X13_3,im_X13_3,re_X13_4,im_X13_4);
fft_radix5 FFT4(clk,re_x_6,re_x_16,re_x_26,re_x_36,re_x_46,im_x_6,im_x_16,im_x_26,im_x_36,im_x_46,re_X14_0,im_X14_0,re_X14_1,im_X14_1,re_X14_2,im_X14_2,re_X14_3,im_X14_3,re_X14_4,im_X14_4);  
fft_radix5 FFT5(clk,re_x_8,re_x_18,re_x_28,re_x_38,re_x_48,im_x_8,im_x_18,im_x_28,im_x_38,im_x_48,re_X15_0,im_X15_0,re_X15_1,im_X15_1,re_X15_2,im_X15_2,re_X15_3,im_X15_3,re_X15_4,im_X15_4);  ///////STAGE1
fft_radix5 FFT6(clk,re_x_1,re_x_11,re_x_21,re_x_31,re_x_41,im_x_1,im_x_11,im_x_21,im_x_31,im_x_41,re_X21_0,im_X21_0,re_X21_1,im_X21_1,re_X21_2,im_X21_2,re_X21_3,im_X21_3,re_X21_4,im_X21_4);
fft_radix5 FFT7(clk,re_x_3,re_x_13,re_x_23,re_x_33,re_x_43,im_x_3,im_x_13,im_x_23,im_x_33,im_x_43,re_X22_0,im_X22_0,re_X22_1,im_X22_1,re_X22_2,im_X22_2,re_X22_3,im_X22_3,re_X22_4,im_X22_4);
fft_radix5 FFT8(clk,re_x_5,re_x_15,re_x_25,re_x_35,re_x_45,im_x_5,im_x_15,im_x_25,im_x_35,im_x_45,re_X23_0,im_X23_0,re_X23_1,im_X23_1,re_X23_2,im_X23_2,re_X23_3,im_X23_3,re_X23_4,im_X23_4);
fft_radix5 FFT9(clk,re_x_7,re_x_17,re_x_27,re_x_37,re_x_47,im_x_7,im_x_17,im_x_27,im_x_37,im_x_47,re_X24_0,im_X24_0,re_X24_1,im_X24_1,re_X24_2,im_X24_2,re_X24_3,im_X24_3,re_X24_4,im_X24_4);
fft_radix5 FFT10(clk,re_x_9,re_x_19,re_x_29,re_x_39,re_x_49,im_x_9,im_x_19,im_x_29,im_x_39,im_x_49,re_X25_0,im_X25_0,re_X25_1,im_X25_1,re_X25_2,im_X25_2,re_X25_3,im_X25_3,re_X25_4,im_X25_4);

always@ (re_X21_2)
 begin
 re_X21_2_fractional = (re_X21_2*(2.0**-12));
end

always@ (re_X22_2)
 begin
 re_X22_2_fractional = (re_X22_2*(2.0**-12));
end

always@ (re_X23_2)
 begin
 re_X23_2_fractional = (re_X23_2*(2.0**-12));
end

always@ (re_X24_2)
 begin
 re_X24_2_fractional = (re_X24_2*(2.0**-12));
end

always@ (re_X25_2)
 begin
 re_X25_2_fractional = (re_X25_2*(2.0**-12));
end

always@ (im_X21_2)
 begin
 im_X21_2_fractional = (im_X21_2*(2.0**-12));
end

always@ (im_X22_2)
 begin
 im_X22_2_fractional = (im_X22_2*(2.0**-12));
end

always@ (im_X23_2)
 begin
 im_X23_2_fractional = (im_X23_2*(2.0**-12));
end

always@ (im_X24_2)
 begin
 im_X24_2_fractional = (im_X24_2*(2.0**-12));
end

always@ (im_X25_2)
 begin
 im_X25_2_fractional = (im_X25_2*(2.0**-12));
end




/////////////////////RADIX-5(2)////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


radix_5_stage_2 FFT11(clk,re_X11_0,im_X11_0,re_X11_1,im_X11_1,re_X11_2,im_X11_2,re_X11_3,im_X11_3,re_X11_4,im_X11_4,re_X12_0,im_X12_0,re_X12_1,im_X12_1,re_X12_2,im_X12_2,re_X12_3,im_X12_3,
re_X12_4,im_X12_4,re_X13_0,im_X13_0,re_X13_1,im_X13_1,re_X13_2,im_X13_2,re_X13_3,im_X13_3,re_X13_4,im_X13_4,re_X14_0,im_X14_0,re_X14_1,im_X14_1,re_X14_2,im_X14_2,re_X14_3,im_X14_3,
re_X14_4,im_X14_4,re_X15_0,im_X15_0,re_X15_1,im_X15_1,re_X15_2,im_X15_2,re_X15_3,im_X15_3,re_X15_4,im_X15_4,re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,
re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,
re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24);



radix_5_stage_2 FFT12(clk,re_X21_0,im_X21_0,re_X21_1,im_X21_1,re_X21_2,im_X21_2,re_X21_3,im_X21_3,re_X21_4,im_X21_4,re_X22_0,im_X22_0,re_X22_1,im_X22_1,re_X22_2,im_X22_2,re_X22_3,im_X22_3,
re_X22_4,im_X22_4,re_X23_0,im_X23_0,re_X23_1,im_X23_1,re_X23_2,im_X23_2,re_X23_3,im_X23_3,re_X23_4,im_X23_4,re_X24_0,im_X24_0,re_X24_1,im_X24_1,re_X24_2,im_X24_2,re_X24_3,im_X24_3,
re_X24_4,im_X24_4,re_X25_0,im_X25_0,re_X25_1,im_X25_1,re_X25_2,im_X25_2,re_X25_3,im_X25_3,re_X25_4,im_X25_4,re_X2_0,im_X2_0,re_X2_1,im_X2_1,re_X2_2,im_X2_2,re_X2_3,im_X2_3,re_X2_4,im_X2_4,
re_X2_5,im_X2_5,re_X2_6,im_X2_6,re_X2_7,im_X2_7,re_X2_8,im_X2_8,re_X2_9,im_X2_9,re_X2_10,im_X2_10,re_X2_11,im_X2_11,re_X2_12,im_X2_12,re_X2_13,im_X2_13,re_X2_14,im_X2_14,re_X2_15,im_X2_15,
re_X2_16,im_X2_16,re_X2_17,im_X2_17,re_X2_18,im_X2_18,re_X2_19,im_X2_19,re_X2_20,im_X2_20,re_X2_21,im_X2_21,re_X2_22,im_X2_22,re_X2_23,im_X2_23,re_X2_24,im_X2_24);

always@ (re_X1_2)
 begin
 re_X1_2_fractional = (re_X1_2*(2.0**-10));
end

always@ (re_X2_2)
 begin
 re_X2_2_fractional = (re_X2_2*(2.0**-10));
end

always@ (im_X2_2)
 begin
 im_X2_2_fractional = (im_X2_2*(2.0**-10));
end

radix_2 FFT13(clk,re_X1_0,im_X1_0,re_X1_1,im_X1_1,re_X1_2,im_X1_2,re_X1_3,im_X1_3,re_X1_4,im_X1_4,re_X1_5,im_X1_5,re_X1_6,im_X1_6,re_X1_7,im_X1_7,re_X1_8,im_X1_8,re_X1_9,im_X1_9,re_X1_10,
im_X1_10,re_X1_11,im_X1_11,re_X1_12,im_X1_12,re_X1_13,im_X1_13,re_X1_14,im_X1_14,re_X1_15,im_X1_15,re_X1_16,im_X1_16,re_X1_17,im_X1_17,re_X1_18,im_X1_18,re_X1_19,im_X1_19,re_X1_20,im_X1_20,
re_X1_21,im_X1_21,re_X1_22,im_X1_22,re_X1_23,im_X1_23,re_X1_24,im_X1_24,re_X2_0,im_X2_0,re_X2_1,im_X2_1,re_X2_2,im_X2_2,re_X2_3,im_X2_3,re_X2_4,im_X2_4,
re_X2_5,im_X2_5,re_X2_6,im_X2_6,re_X2_7,im_X2_7,re_X2_8,im_X2_8,re_X2_9,im_X2_9,re_X2_10,im_X2_10,re_X2_11,im_X2_11,re_X2_12,im_X2_12,re_X2_13,im_X2_13,re_X2_14,im_X2_14,re_X2_15,im_X2_15,
re_X2_16,im_X2_16,re_X2_17,im_X2_17,re_X2_18,im_X2_18,re_X2_19,im_X2_19,re_X2_20,im_X2_20,re_X2_21,im_X2_21,re_X2_22,im_X2_22,re_X2_23,im_X2_23,re_X2_24,im_X2_24,re_X_0,im_X_0,re_X_1,im_X_1,re_X_2,im_X_2,re_X_3,im_X_3,re_X_4,im_X_4,re_X_5,im_X_5,re_X_6,im_X_6,re_X_7,im_X_7,re_X_8,im_X_8,re_X_9,im_X_9,re_X_10,im_X_10,
re_X_11,im_X_11,re_X_12,im_X_12,re_X_13,im_X_13,re_X_14,im_X_14,re_X_15,im_X_15,re_X_16,im_X_16,re_X_17,im_X_17,re_X_18,im_X_18,re_X_19,im_X_19,re_X_20,im_X_20,re_X_21,im_X_21,
re_X_22,im_X_22,re_X_23,im_X_23,re_X_24,im_X_24,re_X_25,im_X_25,re_X_26,im_X_26,re_X_27,im_X_27,re_X_28,im_X_28,re_X_29,im_X_29,re_X_30,im_X_30,re_X_31,im_X_31,re_X_32,im_X_32,
re_X_33,im_X_33,re_X_34,im_X_34,re_X_35,im_X_35,re_X_36,im_X_36,re_X_37,im_X_37,re_X_38,im_X_38,re_X_39,im_X_39,re_X_40,im_X_40,re_X_41,im_X_41,re_X_42,im_X_42,re_X_43,im_X_43,
re_X_44,im_X_44,re_X_45,im_X_45,re_X_46,im_X_46,re_X_47,im_X_47,re_X_48,im_X_48,re_X_49,im_X_49);


endmodule





